PK   ΄6V ��<�p  ��    cirkitFile.json�ێ%9r-�+B
�-�༓�6G3�`�!�<t7~U'T�Q��������o�#"3����mYdj��@UVn��F�ь4����������4=����ˇǏ�~T���?tO㟺���}���>=>��S��������ͧ�yj������΃��{�>���ѴMo�����Ks�zh�w?����#(6B������_��������t��an��5m�t�06&��Cc�tx����[�\����9p����Eh<��};��ΙQ�MtA5��U��)9ecM
�!1�9��G��m��!�F�}fCd �7���F�����y�>�Dx�����ç�o��Tr�7ڊo����n/��O�Y]�[���l�̂o�����*>Df�7�l�̂o��ٵ��p6Df���l�̂k4"���]6Dfa����L�oͷ�l�̂o����Yl����p6Df���l�̂o��9���p6Df���l�̂o���`Ńo��wfCd|�ˆ�,<s>3��|�q�'�|f�����a6Df���l�̂o�����a6Df���l�̂�f�s|Y��|Ά�, ��|n�6��Y�}g6Df���l��"2�3����p˷��e���Xh\���"]ǟJ*aCd|���Y�6Df����`#�?8�t���,��"���l�̂o�����l����l|�����"M��j�j�o�Wm���7�����<��;��!!��9Ȓȁ��e�9���`"r�"��9psq����8D\��(�ȁ�p�PC��E8L�!r�"'�P��RL%�Ve�PY��Q��^%�PY�-�Q
��fe�PY��Q
��ne�PY�-�Q
��ve�P�+��<�B�� �� G�o;��P�,���(s�ʂo;�2G�,���(��ʂo;��?�,���(��ʂo;��?�,���(���m�Q���vePY �t@�η�G�T��k��'Cm��.�-�r}�6�غ܂�[`���c2C2�a7ێ� ���O}!s �KQ���q��Be�7�GI'T|��tB]�����*��?J�������*�2��9ʏ�N�-؝:(�w7��� ��a��Z�4�G�/�����*��?�W�������*��?J�n����Q����%�PY�2��i}j�S�۝:(�w��$�����^"s@ޣ\j���?G�.T|���Be�7�G�.T|���Be�7�G�.�]h��?�u����v��q���������hRc��M������I�y��K��}��	�0ۆJ��p�mC����l"Vv�0"�W���`.&r�"f�98րR�u��C��E8L�!r�"<'�|S�v0i)L�D\��<!�Jl��7��2Nm�8J����G	BT�[[���"*�Tq�_De��xIQ�I�����ǐJ�8%��+S3Ge�G	���\��;�[=c�������
5(l-����a{Na{n�nkV����S�\�;[�$5���wqj�����5a1��J&-��4��4�a���y����2�nOP+w�)Pv
�.G�X�Y����]�లsX�A�),���ce籲��SXv�C��.`ee���r�C�[H�jdz+�U�`p�'��&����]YzG� �O���EC��С���[�	߉��hܸ=����� ��7
�`�)0��L�8���S`~e�,?p���wy���L�mZYC�&a��~���qgp���Q���+�����KX~
̯�p�2a�)0�r6�����_�* �8h��S`~�X~��O���J`���,?淾��k�g|K"~pЄ�W�o��4a�)0�R6,?p����J��������+�Z���/X~
̯���`�)0�R��_���_)��8|��S`~�$X~���O���bJ`�����Yi��ŀ7m8���S`~�X~���O���֟���`g�>7�Lwl��F���/�`�)0�Rj,?p�����J�4�������+�ݰ����O����t`���,?�WJ��_�����ĉ��&�sj������7�OQGU?{�[fL�#=8�Y�,*��°M+��G��A�M4��Rd�4a��j�`��7m���_�S	�8���S`~��eyA����i�<D��ɂ�&,?�w{/�<)�����`��6��8�r���O���:�`��c.,?�W��������m]�������+%���C�3@4 G?�8p����J�f��V���B��]7Zk�F�X릦sS�h߷jr�tdR঩��1EE��@���-�փ�&,�R����	�O���R�X�y�N���+E���;(�v��whLف#(d[גc��Aц-�C�q��1`[ג�q;l+񺀃��_fj汷�o�.534�	���M���8L��L]�d߽"1�u���PMl=�ǨF����P/�&��z0D7 ���h�z�.���3��F�O��`�c���U��(;zQ�rX�QW����aeeG� Z�����(��$�쨫Y�;������W��C�ʎ^A��X�R=BvPv�2���R������������0��(�_�aX~e@/�A䇎����ʀ�� ���Im/8� �ɤ�f`�U���8����y"?p���WQ��D~��˯���<���a�_EE�x��C,����� ��X~5/�A����_EE�x���,����� ��X~5/�A��?���*j�� ��X~%1/�A��?��*Jb^���`�U�ļ��8���(�y"?p���WQ�D~��˯�$�<H�8���(�y"?p���WQ�D~��˯�$�<���iV���\r�D~��˯�$�<�����_EI�x�	���-�I ���KN^���/8|��(�y"?p���WQ�D~��˯�$�<H�48|��(�y"?p���WQ�D~��˯���<�����_Eq�x��O���r��x|���޷K ���kG^���/8|��my"?p���U���8|��(Ny"?p���WQ���"8|��.y"?p���WQ]�D~��˯���<�����_Eu�x|�����@ �}P}R}T}V���?^����`�U����8|��۪0�Ã��`�U�����8|��(yR.�`�U�����8|��;.���Z��r}�6�ؖ[�R�t6L��_�1�!���*у#�5�MQ�q��A�CU�E5ccb��1�0���6'�����%��+�����n���ޟ�fPq\*w� ��ߣrQ�T�#�����o��]qG&sh*��T���,�}�|�3�g*�bj�JL���?͝�������ΜL�4Sq��v�Ok֧�Χ]�93f�]P�m{����fJN�G�B(6����2�ܖ3Ǜf�7�o�9��c�7�7�Hr8N��Ta�S��U|�6
����cX�����G(8��-��>���9d-7~b�h�9�,s�Y��f�S�eN�9e8�1�,�㘪��:�`8��;��;��;��;��;���vo��0�~MjlR����6S7;�8ϱ]J���G��������U	�R~�7�&�ۮ����hl�����7C�%oR\���R��Dҧy���H����^@F�4+�LCᙆ�'��g�Z�s
I�f�Á����Na`N��9=���Zv�)���Ӟ�1��M��ƹN7v�*�T��*�]�Zmfey�*���ęI��l�sfI�2�>�9�f-]D�|�R�Ț�Y>Xܷ�i��ݺ���v3>����i������=5%:~�V���5R�
��{^#��g|:�Z�gH[��!�Ms��*�MΧ��&�ӷc�>���H.�
7!��4�6���*ׅ�i��6ҧ������?��}�����Nz}��'�����^�,�]ݹ�`�K]iw�a�.0ǘ�W�o�Gϴ���G�y:s���u~���c�5Y�����C��N1��<빺V�Ce��!Ia���NB�ڶm�cM�އ�?�!;"m<�۔��Շ@��	���J&
�d�� ��Б�xݱ>� ����V��=E\��a ��qZ��S���n ��s����כ�wz�gM������8�����KLz}��^ߟ�I��{�}ߍc�\�G�56�s�ϡk�I͓V�s�(z �������0�Ly�}&?���s6��rS?�����י_ߗ|HiHc7gߡ,���4]t㦬˓��>�'�~0�S^g��Wet���ƒˤ�^�)k]v}��W�4����~��g�˳�0�!w�Ӥ~j���sz8�:�����~�˲ҳ�^_��l
�<�l��7ַG�Nz}��*�co'�x]\��Mo�kb釔�a�_�?n�R�]G��ɾ���>��);��nmj���G�٘���h5����6v}�ͨU����Q��-p2֥������׵u}?�6�КP|�qlZc�����X ����6��F�ݽ<=g�9��}o|�F5�lZs$r�v��̯��.�^Gׄn*^���PO��u���h�W�(�����w��ϣ�?�L��F=g�{�����Γ^�'Oz�`�rfrw�\K{oS�vb�g��OX2���H�˪p��� F������kw�m��s�8��l��yԓ�����%��v�����^���|�(�೼۾��1�{3Ǧ��dlR���&�����^�o;����G7���J)�)����!~��>���#�Ez���g������k��;�g���JG=��(� �~�+�V9)�{V��d��t�3��|���������ӻ��Y�ϒx����w�)ТXF �e�}����+x�4��A����b��ڲ��aj����l�e�>����cP�"JF ��l�b���e�d"qVg�av[-��o��	f��t���e#��>O�c�=��|��ڥ��̂+��U0�v�D���
f�QH�R1�	��.U8@�p�7��*R�Tq��qmQ�y�f�QH�R��iAJ��'����(�v�p���f�QH�R���츁�qR�T�q­���R`v���qR���q��q�bǃcs���f�QH�R��	f�̎��ڥ�hf�-̎����e�pM2LN0;nav��.�@�`v���8
�]�2�8�츅�qR�����wf�-̎?#un�Gf,�Z�_�`v���8
�]jj�8�츃�qR��q��n�7av���8
��ȁq��q��QH�Rd�	�{�?�Bj�jn N0;�av��D�*� Q򊈌��Mdj	�@DF�^;�2���(F�&5I��|��&��O�ԛ8P�ΧJ"#%���D�+"2��&g�qff�	�@TN0�M��r��nB^��z����`���D����l *'�'dQ9��8!��	f�	�@T�f�	�@TN8����8!��	f�	�@TN0;N��r��qB^�̎����`v��D���l *'�'dQ�q�'dQ9��8!��	���[J��qB6���4�Rą�	f�_��9D&'�'d(Q9��8
��WD���l *'�'dQ1av��D���l *'�'d�/������S��nQ�)���TN0;��ķ��l *'�?N��r��qB6�̎򊨜`v��D����qB6�̎�������t��yR*'�F��Kl9���+�f����`�*�l *'�'dQ9��8!��	f�	�@TN0;N��n���8!��	f�Q�@��"�eg穽$ J^�vP%���$lJ^������=���,Ndt>���(yEDF��)"��ɒ�D�+"2}�+�ۣ����|�$2��&g�_��r�29��6!��	f�	�@TNe��@TN0�M��r!}�+��g�u��_KrWm|��,�RM��6��%�6���P���\��\�\r��ʗ����D��M�|	�}��D��FD�VD�\�����Չ�U���cL�z�JpU"\s�,"� "W	�J����U�WE��
F�5��k��W%µ���2�[%ö�!��V(�`�dؖ�0C�$������L�d�/�J�mY����L&�Vɰ-k�2����6�B��d�0%�)�HL���fX��	ƔL4&�Vɰ-g�ed+���U2l��f��De"l��rF[fcA&.a�dؖ��2����D�*��̼�le�2�J�m9�/#[��L���a[j��'h��l�-)[��L��e"l��RSBF�2q�[%ö�Ɛ��L\&�Vɰ-5>dd+���U2lK����e"l��RsE&1I&.a�dؖ�12����D�*����le�2�J�m��##[�lE�tE�������L���a[j+��V&.a�dؖQ2��؁R2l�6[�d�2#���U2lK�.���e"l��R{LF�2q�[%ö�P�����D�*����le�2�J�m�i'#[��L���f�ϫ�2q����6�"��Dؖ�2�:I&t�L&.�2q����D�*��棌le��D�*��v��le�2�J�m��)��`e��hX�le�2+���U2lKMT�:�*J���f�L\�d�2�J�m�Q+#[��L���a[j���V&.a�dؖ��2����D�*�����l��|����˜L\�d�2�J�m�E-#ۭH����e�lB��˜L\�����L\�d�2�J�m�q."[/�_&�Vɰ-��ed+Q�PɰU2lK�y{�e�2���-��e=�zT�o�4��@�V�zT�\%�*�[�W�*1��j��V�^�ޑ(�����[E�U�ku��zT�\%�V�^��!$"��u�-E"r��Z]{�(W	�յW��\�G�U�ku�U�*7�Q�r��Z]{�(�ʅ�zT�\%�V�^�z�AL}�U�/r�����z)[��K��f�U4,R�l�k�R� |�V3�
A&�a[_{�,R�2!���ګ`���	�D���^� ���L(&¶���X�le�1���W/�"e+������z)[��L�m}���ȝ��L�m}���H���e"l�k�^�E�V&.a[_{�,R�2q���ګhX�le�2���W/�"e+������z)[��L�m}���H���e"l�k�^�E�V&.a[_{�,R�2q���ګ`��I2q���ګ`�����D���^� ���L\&¶���X�l��e��j�`�����D���^� ���L\&¶���X`ƽ��ګT!��e��L�B���D���^� ���L\&¶���X�le�2���W/�"O6��e"l�k�^�E�V&.a[_{�,R�2q���ګ`�����D���^� ����Q2������X`� ¶��*U2qYm5S�d�2���W/�"e+���ݬ���E�V&.a[_{�,R�2q���ګ`�'�e�2���W/�"e+������z)[��L�m}���H���e"l�k�^��"l�k�R� T�C�ʇP�������X�le�2���W/�"e+���ݬ���E�V&.a[_{�,R�2q���ګ`���d�2���W/�"e+������z)[��l��7><���Ǐ��O&�Џ���kھ�alLLs7��^?���*QECP�n�X%�������\"%��e���)/F{F}F���8���`tXa�X%���h��`�k��E�äG��Ћ�v�f��y��<q`�3L�|��`�Xc��`��`�؀\	����N#c���[<σ���g���*̢�StS���E�C��90-�-� ��QX�[�[�Ga1��bl���b�h��8��a��-Z��_X�w-v-v-v-v-v-�/Z�\�<�E��q4�p`��<5��3�y��f�M0�Y��<�<Q���yv�ؿ���v,c��c��/Z�M�Yuy��8����(��G0�8`lq�����hqRc;������eŚ������1�� �m�f��.�`Y0�'�)r`N�x�����o�����jh��|3t]�&��t��z��)&���&�P���BB9�%��IBqg�GB�g> 	%���6?��95�X��n�j�S��:����{ݞ���P��2	E��9۹!�س=�uΌ�m���m����L�)cv7C8�.	E�-J�PN�~���OB9��I(���r:�PNg}J<�]�2�����q��=[���z�4��>���o�Q�𼻖2��v`��i|M~�m�cM�3��?�!O
m$X
�i?k{��q�Ӎ��m��Lcc�ũ�fV��˾`H(�l�P���g׍6��Ҙ�Y릦sS�h߷jr�t<o	�E$}�"GB1g!)	Ş�ǑP���	ş�꽙|��q�d-���t]���r>�����	�t�PN�	�t���n{�=ꮱ���~]3Oj����S/��r*����0�܎a��E��==�!ީ��3tJ�s.$��>
)i��<	����`���qS��Is��[DB9��L�N�N݇�e�fk]��tӫ>e���$�l���\.$�S��Y[;�f琣�Ӥ~j���sz8�BB9����.�S�>;ɇ��)4󠳩˯�-A_H(�\T���N��̫����Č�)��ԟύ$�ӹQ}2*��t�_Z��d�̎L73Y�"Yʹ�t}�ͨU�u�sk�!�ݔ��T4��=A_((�\�u}?e��=Mk���q���ث��.t��rʥ�/�ѹ��Gc�M�ߤQ�6[��g�BB�p9(\T���	�T��\�zz�M�S7��EK��)(�1�E�����h��O��k�Q��k�g?��@G$���Pη+�<���mڱ-k9�϶.L�OSc2C2�-�<��Z
��	eiQt���5�tEH�A����~�v7�&�1�̣���|���,��JQPN{��r�y�<���g��}F�1!3Ǧ��dlR�	V��r*ʩ\H(�r�n���R*s@76IC�z}���@B9ח�e#mb3v1�SrO�<r(��Q��%�$���>�i�:;	},�B���q��.��sH�E_�VqH(꫕�_`>=>���4����_`������i|p!�}iTT�{�6Y�e�v����G�%���8�����k~�@
��F ������az��0�����]V� �@@�3aj�]#P��@��������Ym�ن�m3�(��y�	�	f��x�����/'��V0�Bj���a8�l��qR�| �	f�5̎���磂N8���츆�qR�|"�	f�5̎���糚N0;�av��>�"�p��q��(���|+&��q��(����-�n%����f�QH��c'�70;�Bj��>c8�츁�qR�|(�	f�-̎������N0;nav��>d�p­���av���8
�}>�����f�QH�s%'��0;�Bj�k`�~`v���8
�}������f�QH�s]'��&n{f�̎�����N0;�`v��>��p��q��(���d�̎{�' ���X�D�+"2Q򊈌`�v>eR��E1:�0��Y��O��2�(F�%��4���TId����(yEDF  R^�D�6�l��6!��	f�	�@TN0�M��r�YoB6��~����`��D���l *'�'dQ9��8!��X��8!��	��p�'dQ9��8!��	f�	�@TN0;N��r��qB6�̎����`v��D���l j8��l *'�'dQ9�VRpK)0;N��r��qB6�̎����`v��D���l *'�'dQ9��8!���	��l *'�'dQ9��8!��	�&�[��qB6�̎����`v��D���l *'�'dQ9��8!�����l *'�'dQ9��8!��	f�	�@TN��M��&̎����`v��D���l *'�'dQ9��8!��a��l *'�Ge��?L����R=4���qh����T��ؒ�H@��""�sq��(yEDF�^;�2��@@��""#%���D�+"2Q򊈌@@��""#%���D�+��H��ƙm��&dQ9�,7!��	f�	�@TN0�M��r��oB6���Ϗ������O�\����ǟ����-��� ���0�J���Z�HB�JD�\���K��U��U���#��JpU"\s\#"W+"W	�J�k��D��D�*�U�p�1��\��\%�*�9R�k��W%�5��"r�"r��D��ID�ID�\�ײ�"�D\"l�۲�$#[��K(쒉��L�d"/�J�mYӓ��L�%�Vɰ-k�2����D�*�e�UF�2Q�[%ö���V&a�dؖ��2����D�*��L��le"2�J�m9�,#[��L���a[�h�l,��e"l��r�\F�2q�[%ö�����Ў�Ж�L\�e�2-���U2lK���e"l��R�AF�2q�[%öԔ���L\&�Vɰ-�1dd+���U2lK����e"l��R�DF�2q�[%ö�\�IL���D�*��v��le�2�J�m��##[��L���a[j���V([Q(]Q&.32q����D�*�����le�2�J�m�%#[��L���a[j]��V&.a�dؖ�]2����D�*�����le�2�J�m��&"[+���U2lK-8���e"l��R�NF�2q�[%ö�擑�L\&�Vɰ-5ed+t�L�(�L\fe�2+���U2lK�G���e"l��R�RF�2q�[%ö�����L\&�Vɰ-�Ded+���U2lKMT�:��L���a[j���V&.a�dؖ�2����D�*��֮�le�2�J�m�,#[��L���a[j��V�ʇP������eN&.a�dؖZ�2����D�*�����le�2�J�m�.#[��L���a[j������e"l��R�]F�2q�[%öԜ���L\&�VU�%��d��0�յW�Q�r�`��@�JpU"\�k�֣�*����*��D�V�wPoa����ګ��@�Jp���J�CHD����[�D�*����j=*P�\�k�%P��Q�
����ګD	T.nԣ�*����*Q���@�Jp���J��e��j�T^&�a[_{�,R�Ba�L�U[��,R�2����ګ`���	�D���^� ���L&¶���X�le�0���W/�"e+������z)[�pL�m}���H�ʄd"l�k�^�E�V&,a[_{�,rgA&.a[_{�,R�2q���ګ`������j��^�E�V&.a[_{�,R�2q���ګ`�����D���^� ���L\&¶���X�le�2���W/�"e+������z)[��L�m}�����$��L�m}���H���e"l�k�^�E�V&.a[_{�,R�B�2qYm5��H���e"l�k�^�E�V&.a[_{�,R�2q���ګ`�����D���^� ���L\&¶���X�le�2���W/�"O6��e"l�k�^�E�V&.a[_{�,R�2q���ګ`�����D���^� ����Q2������X�le�2���W/�"e+������z)[��L�m}���H���e"l�k�^�E�V&.a[_{�,�d�L\&¶���X�le�2���W/�"e+������z)[��L�m}���H���e"l�k�^�E�V�̇L\V[��,R�2q���ګ`�����D���^� ���L\&¶���X�le�2���W/�"++��e"l�k�^�E�V&.a[_{�,R�2q����ǟ?N?=��C?s3�vh�i����11��b{��BPECP�BP�CP%BPF�@ʋ�^�Q_��_�Q`��`�Qa��a�Qb��b��b��-�-�-�-�-�-�-�-6-6-6 W���������������������c��b��b��b��b��b��a��a��a��a�؁;�;�;�;�;�{�{�{�{�{�{��F�=F�=F�=F�F�F�F�F�F�F�h������������������T�'�ۮ����hl�����7C�%oRoMן��PN���r�M$��^"��v	�G����rjg��\���xc]V�)��Om�먢�g�u{�/$�S}!���	�T_H(���ΙQ�MtA5��U��)9ecM
�\�$�S�PN�KB9�.	#���HB9�$���HB9��I(�s>M�@ʋ����5F�w�h0�<;m|�k۶�v�M41�6���<)��`e((����M��ƹN7v��Ij2��}�V�Y�s.$�S�ѳ�F��ui��uSӹ�k��[5��� ]�i�H(����� ��� ʩ���;=���&kI�Ǧ���g�����t��$�Ӟ&���4	崧���^�F��kl�禟C�̓�'�f���!�����9�v��-�T��9�N����NiE�o((.�}R���y0)���4]t㦬Փ�<,&��bRP0-:�:et�e��u�w�M���uw�S4�j��\.$�S��Y[;�f琣�Ӥ~j���sz8�BB9����.�S�>;ɇ��)4󠳩�sw��r�E�y����˼:���MpM�X���8L���9��OF垞���KkS�L�ّ�fc&�;B$KB9ח���u�ʶ�5]���L����&ȅ�r�3X��Sl��Ӵ&�MǱi]��{�AwI(�~~1���v�<�5h���&�j�ْf?� 
��y@��utM覲l���Slz��9�.ZR�OA9��((�-�|�'�G�~���\Ӎz�^�<�9�3�8"�����r������mӎmY�I}�uaj|����!XL��j1Ӣs���o?�1������x3�zR��}O��H(.�崏|�|��L�>�Ę���c��a26�֍+EB9�	�T.$�S�D7��uI)�9����!]��>��Y�e �P"�l�Ml�.f�a�C�i��B%�8�q��8��r>�=�^g'���Sh�<=������Sf{
��\��}��~zz|z�0����w��4����Oݐ�����ݏ���o~u�$�!�S�����'�4e��u�W~���ِ<ܝ�z�����{�r�Ŭ`�1s!�}ђ>�2�L�d�-��L��>:���PSh�G���շ�-��v���*�zjlU��j_�0��M�ok&㲏Z������0M))�*�ea�ߺL?SJ�p<n���	HE1�X��诩�OS7����H�V�~��Tz�Y\���~����z�t4���X������y֧-s|�/�e%S"�b�mp�o�Xj��ۚ�nf�sF`Լo[μP�rrM�c����g;Ҡ�#ٖF�Cȑc�)�ޔ���5����X���n�]i�X�7�`��mQgV����w �4����g�?q��@�U�z��}��T<�����q�Ď��q������^�b}����;`��vF�[֧-��<�s����p���<�N�#ϵ�K����Pًv�T�����C3���+ݹt8V���oV,��k��� �h�o"Ö�f.kTM�k��"�N�cٍu�f&��lA}��9����
�}(ˤs��k�[_tŤc�t��j�ɝ1����������a��]7�x���#}�7�r���aR����C��uC�.O�2>mٞ��:��t�����s���xڗ���2A}����H���v�3Mf�G�ܬ�*�$���Rű��܉�Q>�ae֘�z���Ч�̣���r��M�����S�s��r,�t3��;��z��z�T�\E������
�xh��>�h���5�ʑ'�֝��x����؛�I�#�MV��%�i�ֳ�TX+��ƐX� �����13�M���݄��׋r&Jϣ�h���&*�������'Y�7��(�6k���h�D,�£qRaE��!�4�ӻ���v��x��'<b	��X�����n�M��#���&�:�ě�:�ɑO��?�!����/����@<	����J��	�u䅗��29<�sB��4�7YX<�Uy�Un��5�O<w�$ �{R�R:�#5{}s�8�s7,8��.tNbtή�B�V`l��/��7T_g.?2��K��m�]��e(��ODYb /a�L]�\Dl�,P����qX ���,|QJs8��"� ��ɾ)-̃�
�S�i�w���Ӗ�!� '�$�[s"��s1�����$�uzL�x��Dt��g(�C�?+1i����n���!�f<�|(C�Z��o(����B`��ص�Vh�*L����"��ݖI�z����&_j7�M:ߌΦ���<��l[%�=�grd�Hh��%�l��H���!ұ�qD:no*&�qGSq=ɿ&6�8ȉh����JbMZ�ݝ������JH�������b���e}}K�X�������p\'sPW�ؓ�=�^Q՘�zg��z�����7��^����Ú�o�⷟�:�ar�86>��9R�#m3u�������A�V�����x#��>	���}�8v��@2{���a*����5w8H���s��B,����B��s������<~�Z�i���L�C�q�*��̓�g+Y/���� �l�1��z<D��E�2�%�f�/)��𫜨oQY"3����Hb�{�軓��o�i���b����g(��J���"Is��������`H�o��B_:�Wu��|�+���7 L"�B %� 
��	 �� (p/+ P �Y@�y���.��=6��XvoW	��Ds��$��<�ŷ��u�B\� �q�- �� �7K3���!4 u���}�����B�/���x~��9�����/*ly �� �QP��L�w9���Y�Ӡ�-�U�3�^��g��e�π{�
���>��+|�X n?o�wUܚ�}˛,���my���]��4
�e&�U3�:��^��;��q�k�ۍ.�XCM����%�
pYOv��N!�1���&��}C���"+�}EV�k� � ��XoF2�W)AX�oT:�����J�:��x8���'>#��O|F������@�M�"�E,νT�[�}��[��ovW��\�M��7����o�6��٦��\����.q����"��#w�	or�_�w���c�෺On�/�X2�}x����Z<>��x|�@\��w6�2a�o���7����w�ֈ`�_�E�¯a�������̃��BJ>#��� ;�6?߅<N1x��_�,�7v�e�_�ɂ}}(׺!��!K��L���w�)e���Ū|Y�Wb���p�ӿ�]���%ߦ8���ͷ)΀��P���~~ǀ��:~l�-���aM<s�蕝k�w�vݩ�R����cG��Afbg>��qG�Ox!�z�i(�0B;��7�0B{�I;L����
*�0B�^8�3-�`&N/x�v�o��i�|�,$6#xd2�W����W�B�]9ҩo���f_B�ۢkH��Ot�^ۃ���=/]�sr��ٞ�.Ua��B�$��N
�����ę�)�p}�����]e�"�K�@�^(��/�b� !��=�{���(���B���"X��;!i.��kV��k���T~�,�@��@"9�yI�����8*���̿��C�f�"�6U�y9�Z����]7�к4�TS75���F��U��̠#wW�Ui�Ӊu.#�I���F$�
Sv#��?d�ߦN��8	wv�B�#�Y�>�g�ȝ%Ǔp���٩	V���$�o�6�X�ڼ��;Z���������G�ސ!^?�������w?�׏�T�dՏ���^HO�U��g�'n����'� ���6�?|Gg]2b��+l����-Z'^�h�E)����}9ŋ/$Z�)ЅD>܅b��4����zY�mF�
ot�b�9~�>>C>.�X@������{WK}[F ɰjQ�ӵ;C�Xr3T��+ w���z`��^�� ^����wz3L�W�':+U�,CBN����dm�)j��I8��=P �*F��-����^�cmA�n����7�Ae��)C6�zB�?�!��	�$��$41C�!����^�5��$�Y�Gk�|�jU�5�n_���� 	]{�[��S�/�ER�󡘇�Ԧjg�� �p�r�m�YRz��{�u���]�՜M�Ⱦ���r7;���ۗP�_���Ů���P�]��������	��p��e�╘N��dн"�6�6��o-��L�刺 �1���I��7Q(�������-�}�w7�0���|�ui�`��7�5���R�i�D[�z����&�X��&�oFgS��yM����ОZ�b�$`|s�������6X����-"+�wI/���s����}=*i���B����u.bc�����o�&uF��o�vlK"y�>�S�s�cLfH������ 
��������
��e5�h=��%����'�+e]�B�8A�	(#��m7�°*�����yKҬ
�U�N"�oC�;��6����cj6���7[N	�?�lq�F~�\?���&56)��qh����T��خ�qտj�߈���X-�}-��o�oOd�ٻ�1��|gղ��X���}��,�rh	��i��.�+�>�;�B���tnb�����<c7���c�5YC�G;��?���[���m�7��9�������H�J����w�{�~����˧��������8����~�0���Ϝ�6C?��g�%Q�͂Q�t|���O���0�I�h�� ��p66D9��f��(�Vʺw��H*�IE�h���b9#�7jۊ0� ���ݻ	�J`_���1�Z�|v-bVr�RV�O`t���12��T ��`j�����1����|��"`>�/�6�
��y �+cɁ^�F�����W>F[���<�J�jo7�J`m�����12���c�`m�K9}>��5 k��(�x ��8�|��d��y ̫�0�{9>TZ g� �+�-�(| �j 敏���_n�W0�|��X���1��c���-c����`m-���1�r����Z�y�c,QW��^**-��� k�`�Y֞�Rq��&B�t �b��|��N>��u ���(�
 <{c��1��u ���(�� x ����|���U���m=���c�r(  {����zz�q�B=L�g��h�6����,�&'��>����zP���hb���8�����,�&%"6�q���8ՃȂq��A5[�0� �y��A����yT z��A�����T ;z��A�����T [z��A�����T {z��Au� ��0���"R�==LĠ� ����*�==̼�� ����*�==L��� ���T*�==L��� ���Tj(	����T {z�jA偈�!>���Z��@�o�8V���z=�{Zv��j�% �uB�eU�9I����D*��=LĠ� ��D�
��&bPy ��a����f^�K�s&b��?����MKԊn Z��9E�iPi<��4*��=�ˠ� ���*��=̼�n ��a����f^Ы����ލXTZ [�ֶ��^�F-	��a�Y��NR=�� ��iT �{��A�0��iT �{��A�0��i��R��=LӠ� _~��I�����i���E��:�Z?�q��Ad���q���̪��&X"����H�h.$�`C'������ˬ�w4�I�!��B�,��y!X�r4#IMfDl��4��C�Z��Ȥ���T �{��A�P�62�	 TZ |� B���xI"�Z�-H�mPw�(�Z;����*��m����q�]��,]���m��^u�z�-��X[]����>��������t��7`q��b�)0����g����S`~9t�ρ����r�����O����,� ����ˑ��3�Y���CĹ��Ã�3��1������j��F�6`�
Ͱ�Ġe�`����~��"�<|�Hс
�aYC�%:V3Th�e�-Ct�f���R#Z��e����$>F��(��6�H�q̚�]E�Ё����|	�C0�r-Ct8f����M��!��B3,'O�k���P��S�h��0C�fXN��e��b��a9���!:�3Th���������fM�):����P���h��0C�fX�e�[��a)4��!:l3Th��HZ���P����t�f��Kq
��a��B3,�5�2D�-`�
ͰA��(�C�-��b�q
��B3,�W�2D�)`�
Ͱ��A��d/C������ ̕ :l1��P��=h��0C�fX��e�[��a)���E�-`�
Ͱ�uB���*4�R�
-Ct�f�6�-���Q�EG1k�w`G.���"�����A5�XtPf��K�5�ћ/`�
ͰԋC�ŀ*4�R��Ā3��ZtP�&Ĉ�XtPf��K�A���!z�tT���a��1�C�8`�
ͰT~D��*4�R�-CtPf��KMM��Q��B3,@�2����GG1�8tf��K�U�W1����fJ Ԭ	s%p�(�iV�jք������j��a)���G�Ԁ*4�R�-Ó�_-3 LX	.�OV�Z>FiE	�
��[���� ��+{����S��"]�x������%�W}��)Jw�����rq=<@6�"�VT7�^��]��*/��b�UT7�ǃ�˯��!�������5����nX���_EuCb{�+�x�a�UT7$����P���_E9Cb{�K�x�a�U�3����ࠦ�!�=F�/`�5�/ bd�Y���12�2��_Hm2:�W�6����/� ��!:$3��_x#CtXfXS�� F���̰�B�@���	�aM����C0Ú
� 12D�)`�5
/ b��q
�aM�����0Ú
� 12D�)`�5
/ bd��S��*12D�)`�5%	/ bd��S�kJ^ ����֔$� ��!:N3�)Ix#Ct�fXS�� F��8̰�$�@LF:N3�)Ix#Ct�fXS�� F��8̰�$�@���]�8�^�� F��8̰�$�@��q
�aMI���i�{9�T	��zIB��a�����̰�$�@��a�aMI����0Ú�� 1���̰�$�@��a�aMI����0Ú� 12D�-`�5E/ bd?��[�%�. n��{�h�@G1��T	��z�?j��a�aM����0í�@@��a�aM�����0Ú�� 1��a�aM�����0Ú*� 12D�-`�5U/ bd�[�k�^ �t��*�Q%��b�E���������G�-��~ 12D�-`�5E/ bd�[���12D�-`�5e/ bd�[�k�
^ ĔA�-`�5e/ bd�[��ڈ�ǈŬ�J������~�8}��`��8�͠ڡ���n���4wc�a��C{ϯ�}�|_3�7���J�mb��5\d�ylg��"���j�	�c+/W{W}W��8.��p�Rq�R%��j�f�Q�&j�&�)u������p����pl�+<ͱf��Ś�ņ�ņ�ņ�p�ج�Xqz�pͫ�W��S�qqL\�˖���
�b��v���A�Uj�Uj�vr�N��j��j��:	�k^-׼:�yujm�83��*�3kB����S��S��S��S��S��S�a@YA�Zm��{��9Q�_k��L�~�Bh�0�kGX�ڻv���\��\��kBq46�G�r<���:p]��5́k��4���ϗ3p��zg`���x�q�p��ֆ[s�i�0ܜ��a�Y�=P����뻾i�۫�����uɛ�[�����o$�uw�5��ћ;�K��w&	�>	��6���%����=�����j�_H�o�ˊ;e���mzUT��n�6�H�mo%��V���@�Z�ڝ���������ΙQ�MtA5��U��)9ecM
�H���7dϡs�x��?�;H����L0��������Az�r�؉��8�cKS�����N�;p�i \}Uk��9W�Ў���'"�c����!4.?�X;�&��g��C�D�xhn(�tX��7���:����&��46�]���>+��☝�����L$��̳���u�� .�y��nj:7u��}�&7�A�-�����Xܺ�{��$����SC��ؗ�G$��0���!�m,�����L��s�8k��uzl�.��qvI9Z�MG������$�`EI���}ߍc�\�G�56�s�ϡk�I͓V�s��	"������0��z�}�?�ܝs6�rS?���������?�HiHc7�Y¤�t}Ѝ���Nj��Dqğ���U�����?��>.K-��4��^�)��h�hZ�N�Q�I���׹86�8����0�&�S�������I�|?�C�]��}��MgSh�Agk�O��?����0���|�u�-34�	���R�ik��섷$��Y}g*QC��ʽ;�}�֦&�<Ĳ����LVw��-��#���8�Q7>�l�Z�5���c�d*����P;(�|_[��S�d�ّ�&�{�Ǳi]��{�¡v��?�~�_I�s��Σ+���oҨf��^��Oz������^Gׄn*�z.�)=��n����$D���P�?����O>'���1������y�s�g
��Oz��?���͌.���o�vlˊK�u
S���ǘ̐�ٰ.vow��vT�ު4n�F۽�
����=��:8�6~�c6��71��f��l���%������l����'���<o��g!�}~?�<l��N��I�n<�=���Oz�������d�"�Tlw76IC�[z}���c���Q��.�X���y*����g��nyG=��г&�4�=�^�ɺ�e�n��9��ٱ��oy&{�'$�����ݿ��������!�����?�������
���T�JL_�b���/֤��Q-�{�<��$,���/��!/q��.�G˖ϲ����,{,��Ȳ��M-i���Ʋ)�l%,��ǲ��,�,N�)o,i������-uE�JG��k��������~-6q��K2�A���-���e���7\ycY�^Q�Mץۖ�9_���_��������������������і7By#�7by#�7by#�7by#�w����5sޙ��ϰ�_�,�T�|��*��s�/">_h��_�,�7*�P�*� �E��M)A����Hx�%���G�9o^��7/h?�I�@�����C��2%��Qe^ݜ_(�	�4%$�m-!��%Ozn^�D����(���%�_���yQ�gA<�M���.�/R|�۾"8	��@�ƿz!�ݿ>O��Oe�~xV��I�-򻾟}=�D/F�����bj��&찡f�s��Wl��b�5��N���]T�w�ejc1n0]������+vJ�#n'1ح�k���i9qw��.��nO뉛]��=+����p����f�9lXg
��=�@ܩ���l�'9l8�r��O{�!����}Y�5�=="&Z�ؙ3�gۉɕ�����zn&+ou�fof!�v2d��轙����^�ٛ9����l�Ԟ="楲��lXc�e7zʰ���gܘ�ͭ5쟦n������p=���^��bX��2d�1��=妦2b�-�8t�*{�̡�{.$1��=G5���ɟ��Ȓ֙k�y�Ό�7���ڪ���b9O�`k��Ew]����`k�{���(ct���kF�������2S�]l�y_��eal�`踃�ke�Y��2gԽloꉾ5#Ŕ��<��_ҷ���-+������bR9o�D�o��|��W'���9%�Ľm�k3�g��V�I�(r����Z�e�<�����S��A<��w�j&C�7?\�-�fh�/�$/���3'��Z�H*��gދݳ<��mg�|����x����"d7<P���F�Sd�Z�{�>1��O��M\c�qK�F��S��,����q����{�Rp�aW�h�xy����xa)����^�G{숇��=�v�����Ǳ�dB���������I�y���ڳ���o�ֿ�Z�S����]]&�S��?/�ϒ�⎵3g���P�Ms���lX+�{�t�9�k̡݉�X�6��v'["#VJD�:������~��駒�uG�������_-�w���������[X�VR����ꧥ<A�iY���핊ZSQ�TԚ�R`�ͭ���o�MP�&,����y��m���s_{�ZKe��]~[r��~{��^KL�JL�%�_%��ӯ�����W�z�Ӽ�4k���f�v�*1��y�b6��W.j��k��u��W.z�E�r���ھu��W*k&��Z���A��i_�g�=�k�6����ZST�)�9�����o�I�Y�W�fMӼ�4k��U��Z��k����]�r�kA��6�u�gI��`_�`�m��Zd�Zd_�Ȯ�Ⱦj�]k�}��]�Ž�ŭ��^��6���{�ϹW������of�����k��W���X�k��	��	~����цW��?�9��駇�&��Ǉ�>��̶$G�����<�:=8�~H_�/�%��o�y�i�?�+�`��O]j��%�>�&MN5���s�7_A76��n�Za������hb�������5����X�d�'d��~�%�k���Ӈ�Â@���b�Y�Q�|h��W|��w�l��o�3�r���{�?�|>�z���ݧ.K���_�������Ӈi9G�ǟ?��0�_>=}�X�N?v,�]~}��_��~-���,ï�_?~Ȣ~������w�&��q.,�LO����O��{���_?<��4��`���c��׹>��4=�����<��~��`��� �ç�Y�5������}#?؛�ˢ-l�[�x�l[F�F�c/��c����Q���U��}��˧��������w�Or�u�����sQ�O�O�Ko�V�;f�������V��{�s?|� ���������w���c�W�w�M������m���)��`��n������*����̜շ����x���-'���;}��6ov�_�${k��&�ͧVm�|j%�ͧV��|j%�ͧ��Fo>�֝��ֺ���Zw7[���c뱳�����|,��V#|�)���c�dӱ�K	���P8�@��Y[RӴ��)ZKj��+s���7n�������綿����:ܽm�s�����i��CS����H��;����O�����и�;��~�M��6���4�W�[������^�<��}��^�o���ڷ~lS�֏mj���M�[?��}�Ƕ�o�ئ���Ծ�c�ڷ~lS�֏mi���-�[=�־�/.�?���~?<����˳w�~P?�9�߈pn����obx��~�����5���7��QS?����5vHC����Dk�7�{�w�ߓ�Y����^AJ_�{��y,�;_ۏ�v� l�۽������Ε��a�R��ǯc7?����_������x,}�C�_u�g3_��	e���<ύ�]�ai��)��r�;vc2K-�U'�[��z��2?����-����O���e+��'���[5�oN�Ϗ�к�,��>���h�ײ�}*{��)�@�I�tը�q���J��%������Bޭx�}���2i�(����Z�׿��I����=��~�Ėn�4�c�����X(�m4+ڢ[�x�a�ޗ�_������}�a��������ۻ~����������-�����϶K��gK���?w����{����a����?�"A��Զ!o�l�mq$���?MO�l2���O�����S��K?��e)?�^�*��-���Y�<�g�_�
醙]��������n����}9�w��W,oH���'}mnR��:&uR�}Y��bf��s�7}י�~L��%�fRf�6qp��HR*�	/�	=���|����&/��˪��Ch������BPSk���qݬ���c��mh��ޏ!�e��F��Z!4�+\�}�%RZ�6�w�"����R�?����~�b���٭|������0N�eh_��"��6���y)�v#6Rq�{��n~�.-��q�������9����ճ�����>�o��4��eo�[{���s�����G��X6��1:���Y��֛p�6v���7Sg��gtv ��g�F�-c�*B"Փ�쀄բ����r�1�gQg>7i�i�ɑ�{u��6[��eN��2'�7�B{7	p�hREZ$��}��z����p�̃��U�l�rփ��[�Q�_���>���Z�����zqT����@�&tB����n�B3LJ5ڎ��K���qTq�D�bI�o��'ެ{�x����A��n��Y1+����Y�e�;��H*gJО��ʝ�q㱭ٱl�fǍ��2;����Ռ�3"�p/mF|f�5#�p7�J���Ϣ�9t�2r<�%Ր&��e�v��祘�/�.������iLX��|k�>=vcn��� (�Bv�\��~]N�U���`�֐�(D���s3���8x���ߨ�Z8E5̞����oab�3���y}�+_��M��:����W����3�W�\�Kv�������߼&�����??|��o>{y)�������׏��<����&~!s�̗�������_^������[y}��g�!|9����˯_�n_��������O����±=E�E����<���������#zw��J�<Qyӆ��A���d�۲V�T���ݺ���uv�Sv+T��ώE���u���v^��RJ���^q+��'�����^6�b��{��b	��5I�g�jB�I�fltWr��uM�5�\7�<���Q�E����B��}���Ͳս��+1�.k���\̤�����Km���&�B��ư�I��Ђ��.޺��`�at��/
�}+�U��	�����q��);�\fC�f������_o5�/+��U۹g��*��$�Zcً������LqS���(�`L�3�mt?�����<�:;��41��OC�3el��ɪuN"�N)�;�"����e9�K������W�7 H/ۯ"�/.���t�))fm��l;��T�9��]oy�,gݗTN��@���3!;Ǖ2�b2��_\,��b�p&���>,"3�	)G+!�_�������m��/���k���S��Kp���ܤr���͔��m^/W��m��e�U�q�7��J=�������巶�!�e��Ǣ�*��2���C��U�o�ܕ�V�U}=�Kң�w�%��巗Leg_~Z����fR�A�/���/�Ѵ�O4M���Iw;R4-�}M{��^M�_~�g����[���-A�ʡ�B�Q'�^���fM�ɺ��9��R�xXvBUXi�s�ۭ������'��h�-�`�ߔ�sI^�_����7�X];�sw��%}-�l����/5c�}qϿ�V�ge�`&�C��k��f��D6�a勓���V<O}m��~˟�y���/ۦϊ���]62YٝY�_N$�Sƫ�vm	k��a��e�%�t
K�?L���c�Ъ�H΅^���Od����i���KV��i�����������Uw��]�~���߽����}ҿ{��w�9�>�����6.?]�E�l�8B/O^���?��[��߀�~~����o�OX�������]��w�o������������P���1�����)���$>usF��C�6��������ݿg��՞0�q�j�j�k��j�Eh����/z�.<�ր��Vy�=DԞ�l�y&j�6r���j>ӵ��A}*�UjO)�t�O�7�9�����Za�g�����!j�S+#��a����H;P0���h�;V8�Z�U
7g����r8Ѡ8rw��?�'�7w
л��+����Vvw�)���fw�=�cO��&����� �xqtWpEv����v_���}*�F��S7���O9����� u0�q�G7���.�w��wO�mǢ�W3v�ۂtԧuJ�s��fp�Z�����ЫU����]E�{�l>��t�R�m���sOm����R����Zc`�*t�^�W�B$���)�gݸ�Q$+D{��٪ynu���p�f*Vs*���\Z�I��/�=e7=!��+�m�v�ťiW}|4��Z�qZ�X�<T�^��jY"�^wO�m�J�+��ݥ���TU����]첎���
��e�-��e�*�_���T��/<e����;���}a.�TpE��]����۹��u�p���r����$J燊 ��aN��W��wjvJ6�����mo�6��=ըv��&Qb�mJ>vSD�P�Ei�>B�eEr�VA�V�n}�=
$E�}�I�*�L|��Aq�u/�6�i���4��ï
zL#��}�{S��~�ўj�״�fD�ST=��'iK����XN��ҳK�I��jG�҅����g�v=��U�Z5�3uA�f�s]�:Q7�]Z'��A��MKe����]"=լ«��7iOQ�l�b�foD�.�#+rk����Rn⽥�ֳ�R����o�Y�]�$>Eՠ,tp���um��s�GX��ś�=۞�ԭOEz���b�]�$>Eֳ>F���%:2�-9���R��m=��vF�=E��Η�������N_k�����m~��o��W|�̶A�R���6؃�N��{���ֹy>I��U �`nk�tg�j��m�K�d��F����q���^P��N���:vo�����KӖ�i����jM^���W��T�d��=�}V�&�'=����uV `��$������VPN>��ڻ;�wOQ�a���I�T�|�I�z2�3O���ν�/pϱ�{�:���%h�-�>\M���
��d	�)c��)�9Ͻ�<��gzO�������5����۩O��C�N��S�N@���z=��g��4C�N�_�}�>��o=<bwA�jmSa*���U���Tb�Z%n���T�~�1jJ�<��KNn���Ǩ]?M^��t�,x��R��)�����v�����)��qs��O{
��Y��#_��:����?_3�"_�ʚ��SԸUD,v��֭T\W +p|�|�"-�_[�Q o�)@�\��W*��ŏ{
p�U��}�j8m��t5���=������m��wO�������Ska�pիى5G*U?,�����!�M�"_��o(6��)�
Z?�&���U ���i:?Ë@���K�����v��C{Jm'îb�S�U��ݴ`mo:=�򠺱��MR�ʯ�wqj��sЉ�TS�m7��*��'in4��lۏ��v&#u.Ӟ���WwӟD�+R�!�n:�j�����z]�����=���՘{��=%q�r!�.���Z��Qm��f�IC�����~�G��٨�h�*�R�:�ZŹ�s�����/����I׺�֪��ku��,�W����K�,OU�jyV
��������Z���v]�E��"G[�n�G[d�x�D[/��}�[�]@���o����k��{#�����j������
�=�MU��q�Rt��T�����*��
�=T��f_�+ ��崂��a� �qT{V����s�ؤ^�Wr��"��zt�:P!�;����y�z���1����W�X��p��y��gx�\�Z����5w-�q�0�_�\���{�!����,�i�nz)���졢E{D�i.��$j8C`��eW��pb���d!oWҠ��T�Q�n��Y	�n[������+�.�-� ���XFޮ�z��\	"����w�̆K�;a�Ӱ�@^(�.߉�dQ��&��Cm-�!�(�Q�c�S���}���D�q*�V9�LĻm�?�s�
}��8�5�J�@�`�8�>��EeW�q�%U˶ �IW+yp.Eaq�kWz K�ׅ�և��E��La�qj��h��/^+��Q3�E$�_�av
����{Q�����7).��p�g�?�G\L�n�6�J�oB���X���&>L�I�룒� ah��,�Nu���g ����lՠ�MBx;��׀M�򸦣!�5jI^Ҹ�����0��v��{6]�gƷ�˽�Ǳ��k�8�O���{��ɚ��Ӻ#�̄�h���4�:�ӽ���\��(ەnYs�"-Y$��1�Vs$�&2�v�G�Ь��"y�Й�7D1�f,(*N3kD{���?(�S6ֺ0���%4�zԢcw,:�J#L�u	�����j?WƋ�F������ME6�[��C&|�Rt��#��S�����Y��e��Ɲ>l&�1��"�ɴ�e��
�2��������~Yk��le�!���kߔIvP)�g��j6��bC.�/ue@6��Ʊq����}��z�	.O)�iU��hB��� ��8�QE@6�髶�3��H�<�����8��oJ�	�9&����Tb ��rdfx�bV!;}n�}r�+J�<^rŌ��\O�솹���(@�X�U�ӗSw�^Ǉ���������\<��_.������^��|���o����zz�PK   |��T��� �' /   images/13cec52d-3863-489f-91e2-31075f0cbf82.jpg||XS۶��bl�E�BSz�*�Pꑦ��ҋb�Jo�$4���.]���ti���w����}�d�5�s�1W�>��?B����XC��&b���ڞ�X�\-�< h��������m9QQ���uKs+{�;�o��9+
�W�s����������bu=�����䕳Wn_��is���J�S�`�ig!kɣ��}������V.׹���"9��Q࡟\�������b���o�zE��������Ya��gŸ�eE�IIHH��;+vV����91�sRrg%��Is�~�9YZ���4~_|R�������������s����g�D�Ą���$��w�IΧ��A�����涋���|����E���O���\����u���E���삷����v&xܶ�[9;�:YX��O��K�߇�;����8ـ�\���`�joEr�TS�[D,m,�Ĥdĥ�$e�--̭���H��K�����[�IK��37��s��v�ąsddd$�.Ȩ�;��*+sAVFMLFCBEE嬌ԟc5I�.�IV��������r����88n�A��M���/\�Fؐ,ܝ������������=7}��l����-ωK�K�����>g%qV���������������uqs���[���w 
���g$rb�b��b2�b��2²��l2V���g�YK�=+-m!�#
�(��P��+ M��?5>�SUV$PJN�f����9�,��ɰ=݃���˄`bbB v11�B�F���̻���nf�H$r/�~�� �b�����k��ݻ�33�?|p���(�K+}��?,�,��k�o����ޮ�L�#++��k�b`���?/Fxd{��2�o��s�&��]�,#�h�ݻ��V�]�B�;�[wd�u1�c@D�*>���4��]�Q_?:E������g�|W��ط�n5�3�h)�{�hV0&Į�̻v32ѯ�
.�s��G�;���Pi/Ĝ���UOK|��h~��oO`��� ��	����R�V�goC�4�'�`p�C4c*�DqS��Ac+������	P!0B�,�T��n0�1I ��B<1D� u��֟���Nx�ҥ����/�C�T���(J���*Cg$�� T�|�33��!��Ay��vdC��} ��!����H�M9B�?��'2�£�gNSF���@he4���?��.�@2�B����23
JS��#pqD�<��"T`�9��C�R	��KSQES��H�?+�CQN�b��S#
�p��C�H�2v7�]� �s�?�|���1���*@�NC���t$+6x���¢돢��� ����RA`� ]�=F| wHc*�� 1� x���:�
�Q@�	�F�{H�r�H��F����<x,�@M*���F )�X0�ʴ&1$�F��ʖ�2���MމN�n0� O��� e
�a����	�B�l�(0�d]$8&@��.�	r3@F8G�4zN�<��0<��!<�4�T8�%!ڿc��A0Y����T]����VGS���@�ʙ(�`�;�����SL�! �.�?U�Mf��`Q@����h���@dP ��GR�+��フ1`V�VBz�2�&�"؃�M�/�2�T"3�*����pVFz!�ل ��N�(���B ������R�L(X�.�	'Fon�K�C��>�Kh�;7�I��|T���h�l((�C �B�@��� �ƞF��X��e� �-�{�n����
�B �tH����SuA�R�P0
� .������M撃�����.Ai�H�*`Շ =�ȇ0r8Q�N��q�Ǫ��J������T���� �D=�T�h01 ᥌Yp�u�r3#q0�(DO5�J����OtA��q�!ɂN#����ӓ��a 0��g �݉$��A�~����9���a.��@#��@�h�]�h ,4�E7 ��A5D��g ��
g�!0����颉j`LPE LP�l`x�@������H���(`�D/2z���&���t��m FT��{�D��z�����A5�9U�� ��㌊2
�@�Bj;)P�(��K�����	g���<06Ɵ��	�esKeSP�D��D(U7�3�YL!T�[>�	�xV�iU�0�h����^���p��l�0!1�(�e�p�
���� a��TF�Щx�M (.�2��.�D�;����a:@�]�� �0��@8�#<�� 0m������ �`N��`rAZb�qP���E�
���� �J����0�7�%��1 �KSf��'�`L4�*��ac":��Nf���A@�Нi�2� �a���!���4="��
����>D�`�M�ˆ1u�s\�/�1��.x��AWL�Ap����"X0T ,�L�rؽO,	G��¸� ����g�<r ���HU�ŝ
�@}�͟
s1�	0�F?��4�Ee<� g`�!(��2D���7�g ���$$�.J��;Uop	P�-�� ?�'��Z�.C�c�]6�@5��&��u	���`������o9��� ����T�����;���H,]S�Le��(�ae@�l�������E�'�@݁$1�k�90�.�D8����1���py�A��D�%�L �	s��:DEmg�wp�(5`m����'��$��C`*�8��IP\�m�;�HK`) �;�H�J;��jD�<}�����T�^����?d
rsJE�����#
�oc,R��a����龥�;������� �t$�A��Kt����9,��c��$��0>� 5�A�]�کy"_(�S�t.��H�l$8�K�.�ߙ� ?�tL�JՅ��0K��ǘ���%�'�U��l�� ��`p��#� �?��H�`�A��r )cv�B�iɟ$���]��13&�� Re�#�𠾐H�����.���
	���{W�� xD 4���้�0S�8A��uQ<�*`p���*."����%0�(��_�+�t'�@�wBU g���$H��3�
g��E78 �k=��o��N�1�M�� �-�� ^�MC�
̯�̰@�} :�&��jD z��(���)f�Kg�]l0y�Aw4����DI����]$L}���������Ґ	�� �	�D'/�#X���33PJ�B�z+Fga�Ɏ˂��`���3Âɳ����j�"0t�2�E�(�PY0��`���%r����,��M�=�f(Ɗ�n�����oh��~w)0#�� �;`�AQC4�� $�ς�������;Ђ]#�E�A̩t%d��,���.��?]�.�N����C^����t����SYP�^�D�;�'x61zF����%a�N��)t&�7r#`��E�Y��7P�'x�z�u@H2ʟNˀєw� �^���8v�
�2e�G/v����'�4�-�?@�� z�HK��U��B0DPp3<=��Z��T��(��c~[L���a8@[��%Z��E���];�����!zB># G)3���E*�Y��z��2�[�d�Bҭ�.�P�A�dC1��`6 71���d&c0PY��I��tG�E |���a��ג�[1�d���P
�:B��8�8��1���G޹i�i\ʺpx�8л�Τ�/�>���-3�%T�w�t���&��[�Y��,H�@����Gocᾐ�b&��]�)a�k��9��!�10!<:�L�{G����� k�a F�j��s#�Av�P)�u����
 -H���Iw�,�`���;\���wP" %�Hht�Ar9��L���Ā��7��E��V }��1�������I` �
�I�ENM_�Y���@��L�lb�S��ɂ�TTz#^�Ņy�#=da����ÿ1��b������E�B�-p�ap;���=�jg�J	�uj�%�߾�4� �"ª	���>8S(�q&�М��@OE�hc	�W���4|��X`���#�oѿP�A"`7�X����OZ��(��z��v���N�G�q\i ���!�=d�:�Zh
��vM:���:m�������o��Z�K��X�TF���o ܤ���;�� ���:�6xF���\0��,FЭ<>�����S3#���#��|J����A y�[By�N��:pn66Ќ(�q��q�h ,�����	���̈d��0��!�b膌Jo-��X�U��BV ��>F�*cf��?%�OeP�	�m�O�0�ա�f�,�4[��#Ր�ݜ )�O�p�j�;kF;&8� �	�.�B�p��C�W�`���|��-7�4Hz{Dxn4P )ʴTX���wǧP�S=X���8���~�K_��Sl*�u���w���;��\N��=6m��!0Oi;�4KH /$��:dC����-�C�7\t���	�E��v�;�G�±nC��N���:a]�D_������S�� ����������M����k^����ۢ�>�]3�4�) �x�d
3�K��̿�N����A�`�ӑ��/��, ��
w�H>�Fz���^��5�`NH<t$H:
b/�������җ��"A��/���R���A����C�'�>tX���ow�uz3E 5ۙ��P��)���v8o�ڀ�% ^���i�B��0x�{"� ������`	�p����aË���]�H�3/8;��x���j�5uF��llp@��V&钀�>�>���H[�.UW�`�
�pz*�95���0��Q&���!x�g��`{�a�Ǡ���ʔ�En@�z��Z���Γ
�!��Ѣ���vV`'N���=���{��s�Us^��[�sy	��o�H&F:�3>UW�O6�:X��N��('��娧�S�P�	.�����������l��k�b�����5�D�G�ɵ�9����Д����^Q������͑����R�8۹ϥ�'?Ѩ�:z��{�
R��X���e]��W����"u�M���8k�{=�Ѿ�eѳr(��@_����q
�	�ᦧze�#-��(j�J�,n��n����>�%�nqQg$�]p�^$n�������i���j_7��z#�fL�u��Y���d�~�B��lD��: `���E��I�������5~/�_щ���0;��D�~>���L�Ȉ��w�����}� ��)�&���c����;m�o~�����l^X	�~�h��"<Vc�C,��Y��^_�O��_���'ns3y��^�/�E[���sba[$Q�)��&�;�\�̪���ԓ��ڂ�zO����~)�,_]����ܤ(��^6��(Kq��� r�����f�3K)cl�qU�n�[{ .���|{%mKO��`ъS熳�cNT�SJ4���������wO~�n��nC���WWsW$�F�6��9�yH�mh�E�:��zC%7zF�hZ�����#L�GX&���X�/i�}�#�L�>�}�����h&�xr�4a&��1Ų���b'|�H嫘fԤfw0��p2~-^���L����6VW��+�B-�E��;��Uf���k���dblJ��^qVR��I�w��1�ɭ.16{�p*�lTG�A���3�����m(�PEJ���Uo��<�����)����44��o6�ȝ(���OZX�qސ|v���ׯ�x]
kZj(�ʘ�1齻L-Q�ʦ�j��DB'��LDy�l�}�F��ē�
�ehU�\���:�2YHyܽ�2T�֛P٤ĥ-��Y!�-s�vz7t�/�\Mh��2a����^�j��Ƭ�)�Q�}�KZ����nD���JT�H������NY���Z񍈏B)�
��f�fZy�!j�P��F�t%��v�����ޘ�_+��+E��[��m���eoQ�˼�,����K�;iG����V���QwiָX^8��r��ɺ׳F��-��V�''����^�����Ǜ(9��&0zl;�\�P�r�>������+nF9F�>B��䗕V7N$Ĉ�i��~���{k?���O�z�L���O������tF�b�i�-�̋�ay-����eo����Ji	�KN��>�{�����N����n�}���wɯ9�ez���ߨ%&���LQqn�N�~���t� cHlkw���X�z�uԭ;<K����G�~?ޯ����@�3׆�vߕ�/�J�5��\�h��g�ޅ�Emf�\�f�����6JiX>\����ԁ1���y�6���,l�:��%XU������t�v>V�z��f���6����O��_6&�~�f�n���{Z���w'��a�~2����g�޽��z?=��)ɞŻ��y�0��^���S�Fc�
�)��d�O��#��|��l��R����&j�׹�{���Et���ބ��L=��]\g,�'�4����"���Ù��!�/u��"��c풥n7l~�rl�P��v�J��\����]\����~̦�}+��6�3�@��T���3�%��1�Y�ލ��;:�����&B�+�~���/+7���ӳ\Q�¾茏���ƙ��ڇ�?�k�ژ8��c�)FԉR���l,ۺW&#�����"�KW�V�[k]#�7�k �-5�i��9���o&ݿؼ�|�/'g��S�A�я���J䑞Ǵ��a�
����;o.�Xe�,ğ/��<>rf�X�״���Z�\��Ϻ����E]�+�Q~�"��.Gd7�8bp�i-h��˲A��]X�p^���/�Yu�=bP�������ԡY<8�%d|�Y��[G��b��W��.�~�r��k���O���\�~Q�~\)�~㓯Ը�Hd�p�MSqU@C�:>�"�_;�w��$zz-N��Iِ��G��&��k���a3o����B/�^p���j�;ېՐEѰ[C�:�q����oq��(��T �nfݻ�t����E����9���GB}S��¡3�����WI3��-�=�OKռ�S�vp�S%*P��h��Мԃ�#��7�.�P�ٍr��W����By�Yɦ��o�i�R�Ճ�U��B��,�2ݍ���("6���uw��w�nm]p�η��u!��b��x[�`�X�ρJ�h�؎�=C��^<��������ɂf���^�"�+K}{��.��=(�.��iوI�u��Tx�5�ؠ9�*����s���B/�/k��Q]�F�M>��u��r��y�ޮx!k����B����R��!�f�:�bߖdQ���rJB�]�/5�0o��u��K3���%)�ul6t�۬���K�h/?��w)G���Y�D��{�g���Ӛ(�����
��j�J[�>�ʬ'��I�?�]`�s!���`ن�i��b�Rd�ZI�r����/u�D��6�������t����>��U�K8��7�N�Č�=�y� �|=�p�OU6��������]�f�Bݾv�v�������R��٣+W�.�u��W
�������A�^���'�ېL
��φ�qw���F�JQXǤ���+f�3?l
.O4�|���S�o���b�Gb^�����c���{'��>r�\���1��2�c��F���{}���+ál�#��������fI>��y�)@+�R�ʜ[��W]���H'#lh��=4Ņ�я"]����~|�r���[ش��*��`�t��5�ǡ�]����7�?���7�y�Yf=���v�.��>p�LD�B��𯿤���|/�,���@�k,D��q��f��%�u���&��!����ΕI��v��e�R8da1���L��AuJJ~�����6�U�n9j-e��ad(�Kc��������4��-J?�W|?�j;b*�3�;�����c�ކz$�v�u�$�V#ϛ���s;Z;�"9,�{s>��z��\�K�qe���eB��Z��c�-~��Qm�m�k���K̼�>ԶwL����F�U\ԃ��m(�e-l)k*�������Ht�^��:���'�,6����s���ҋs��z&3��]��X�P����rn`�V�n��64��=��O��,i���L؉ꩆ��Uѥ����'3'�ݪ�h~�a��e��^m-\i�/��~�X���_��J�>�C)h*�l��񏂝��jz �?K�(І�\�	�{ǔWRE��?n8>F��.��_�S��|�4������]�\��O���V&ϧ��>�߆�}YQ��6:����Q��W�z�R���}p��1��&O�,齾�s~��f� #\��5G5�2+��3����N�R+�����c���~���{���'yխ6o(�`��������mH����x9J?�,� �3�<�]tR��_�=�9c"M�؟����� ��K�5ci�d���WM�)[����'&R37�������$B؆gt�yy?G�e0f�J�f�׶�֚= ,�X%��[�چ(fd�0S�M��9�iwH�d��I����+�J��m�ڏ�h�f�ն�ן�eGY��eˢ�̠����Ѿ�5麗3�:*�^���}������w}Zݠ:����	��/~�tv�f�����O?E��*�3���w�V����0Q���38���p���6���i�ѺV�vF�;#��͗kN���X/,�F���ù�G}�����߆KʨΏ�=�~3��&8���2Wf��v+��q�O��v�r���O|v�V�ի�U�V�;�x�X+Z�u�z$_Qbe
��a\���g������£&!rF09|���o��r����,������mU��ߤ�:��_ɶ�)LPz]��ؙܵ)��J�윯��ާ���Jb{���P�h���h���.�M��D�4�bl��b���Sn�mS��Bl-ɠ�=��~�G��F����+4��6�^��z������PmH��"�Y�I�M�ҵ��	QN�e]���[q�[�I
}^j壏F�D��H�nm�qw�Բ�up�T�]�`�=?���j}3Dt���eX���g��l�N*��N������D۠wU��~�����jF����μIɡ�k���9�H��P-�h�q�{��wj�����G�#�]]����黽!3��XF��=<-����
�}��x)E?�!�:!����Q=ǈ�� '��*�T����.��v �j~?�n��p��k!k��DZ���q�	�i��Z�D�X��P��}?ʗ��o�ךV:�O��\��2�����<�6���IX��h�غ�U'p2���ܳ��&N�&���@��п�nZ-�� �:�UZ����[\�&Ϋ�ęK�geA߈���5�X�m���nD�f;�	7䅴V�&���X�"g�r?՛d�5:5y�΅:]��$|?'�T�\�j�G�Qm���m�V����e\9�/h�����dJیתpj૫-~�t�w��z���cɊ��Ļ�P#������y��fx{J䏒�X'ǹI,��b��cX�%M�J���gޙk_�n^n[�4j���{�F7������/ǳ�7��=��KS�?~t]_�鴭�ǥ���&^gn�*��^�Y��[6hr�ۂ����Ί�!��ٯž��^��
��;�'\z>��_!M�DW^��l'N������:48�jm���%vȂk��b��ɵ!��r��9牲	�WC�N/��"'z��`ޜ�cP�wr(~$9Vm��ح���#�GX�x���x<ȷа�����M9!��7�uB�������̰TND�c�uT��񗟴�"�W(�H3�KuMd�gB	���+t��ĦT�7�ODV?ڨ<qk�;�z��FC����SW0nUy��*��o(W���δ�_�S88q���H�Sx!Z@�l�C�NX�n?x�r�W�����{�2޾��.! 4����[����B�ؿ�>h���u�ɗ�#���ʐN��<޼֜��S�[׵���Uv�'���E����vY�S�<����Ȼ�Ӕ��ϷN$%�:5�w|1=Y�*~���e��;n#>��|�ZF�Qqd��+Ym�!��kc���i>^��.�֧�=�@�_����%Z�:���}����`&3�
`���eW�a���jR�
&�F����O�[H�on�}V�qn�ԍ/$n�����X��j_^�_�D��\�Y|��k��u���5��{�t����[s.ղ�f��V<�>�ۖ�hcR�.���N��3�a��U����b�x8�~5f��μW�����5�P�B�+aL����=K'n��=�S�������|9��7[}cޒ�����㍮|�(/(DY_�+�fY�qz;f"]�DӋ��u����j���64|�e��"�cm��D�ڛa˵��G�,���MNf�!�i|�������_n�h*�:r�S������F{�������׹�#�*���w�7�)*KJ��L�v�2����W�Ѷ��^�X��U��#/�tҸ���XNJ(0w,�O(�c=��_4���~.�),���b�o����K7��H���Z���[+�t��=��W��kR��kq���\oB	r7�����;���q���~�9l<la��X�̈�k.?��jzv�	�nI�x���>��Թ����-�i?��z��k'����9l�*�QY޶h4`�n�=14C}om����ٹWG�'qß��dWŷLs�}\u˝�9!xЍԧ�$�&�,���.�d�y�mR��	*����뷉�%���olC�BZ�|/Cx6��Ȝ�Ky>}_עt���|���k��i�G�̦�5���5��
�cG�㷡Ϋ%$%,Q�h֧��X1��RC�ƞ����4|_�d�V�g���A��Q�U�*�N|c��ͧK�՛3���,��"I�.�=�ڞ.%-OR"	v�>��OkOT{S_b
4�m�"��_�Y�59���]�>6lz�v5�v�֍9�q�IId�f����29�L2�);B�]9g��4���O[���L)��s���lQ��eYpG��r �0+eWk:F�Dd6�7O}�Tt�#tW"�o�+Z��w���w!#N��ەQ�.D��eD�ㅆ�q��)�O�9��n�a�ZA�P����m�� �|��z��pIY�2�);�Q1,j.��X�~�G�PI���21��[���ھ�{Vw6��^�QXa�mXp͵7,��N�&��]a�;c�8Z��j�~�,ZF�
'�n�o¢	�86���T�+��^b�ƞqȭ�YZ��j[��� �-�Ѻ��Ֆ�ۜ�$g��mH����f��GN��+D��O���&ѽ}��%7w�sv�(��� Q�VL�ж��h��hR6=�_T�W����f�a?[^��$��>�~	q�'C��z;[���2���� �-��LzFۛG�˱"G�w��vm�J�'7U?���WaN:�m�B��k*]k�Z�>�b�-�^��G����|���U��OC��N��=��&��a�K�pg��c��TF�����lQ��;2w��gGE�X��~�Mp���Ht���%�m:+�U4���۰��(:��:�^;Q�Q:5�>U�f�_�����2�9r�V��6�G貛ĩ�=z7'���g���?�Mn�J����j��gŖ|�j�m\���|�#Vx��-������E!��#�!ru_��p�I�O�X���E����o�z5�~ަA��wn44���Z�B�*_�v-fL�f��I�|��Ԩ�x�>�� ?�v�\�Wk��2�����ې�6T��M$���J¹bGt�Qq�gCY�1�ʫ�i>���6��vk)��օ%V;��Ou�'��m̹�C֩4�w���j(�K�8R��t.�X�ǅ�|R|�v�{��j���l���$cwQnK����6����_�'%�q��܆n~��\i�Xm�����}��DVDK���O��J��z.���	��㒩%��9����f��E��z'�S����`nToA'���V���?w�]Q$.��f�o��͎}�z�Y�]ּ}��\�KP���dT@*_��*;E-]:���%�ѿ��@���dr���}-����a�SɍQ��?'Gpv�x���~g	�~z�0� `���`���U����!��6���~�}$���'̥Z;_�L^��?q`������ϟ��4�m��v]̟���J���dX��e�eWr\�.�|1��s�$U�K�s6������Q{&��F�tu�!YJ>Z�X��Q��*;gv��ȩ�v�-k�3���%���� Y(�m6�}��������3%����RQ��9M���ȝ�;u��i��p&:˄����`��U��S}�z�<�����a�,&��{/le˵ka��߹"��U������s>��9N:��y�3L�Bٰ��ԑ���ON�j9T��͆11��ğjg2R���}EK��p��3=G]����:bq�H2�����ٶ~�T�{׃�	x,K��>�����C�RRV��x/�oE�NL�'p�FK�C����OY�y&Y΁��5�bP@�,�Z�tX�X���`���x,�h-}r������G�h�U�S�HnΒc�$��{�#�"��Nٲ
�����4܍rՑ1$+MSo���ԑ�8�@�.�J@�;zJ��B�1�K��+gb\�v��,{��t&bX�-�pP��ا�F��8.�n弙�\p�K�_��6��$�Cx�a�cz%�B�Њ�ɽ8� �������,��tO�	}at�q�]���D��M���J�Th���$���4�r�~�$��"�˾>c�ä�G����p�X��D���֚�U]�y��o�㱆6c�(�:���~�X�;��]!�v9�7�Q4�^ފ�TMt�1k�ٛ�9X��rUEE�+SRGjc�_#o7\�K{ui�H�����'�2^����}���j���Bi"�Iy�r�݋6o��ͳ{&M-<w�n*�8���Y��,�Ǖ돖z+.1��kA�������D�<;�?ڋv��cKM;��%�?�ݭ�6��ICr�-ג�{58T�t^*�S�z�#t���v"~���nru���MM��c��Gj;��[sA{J(j2'$#ǚg��/ה�D�UV�h�1}C�#&o�\&ƿ�>�>����K��S�<�(��q�v�j@p)o�SW�����y$���������z��KS�Ӓ�}��[�{ا�{�]�yЃ�H�kLR��h��G����b,��9��*�����M�Ly���I�7����Տ��}�]R��L�K.N#�U�p��c��w�棂5��|*��fi�n�ؽ�w�1��-z,k�����9	ŝ8\��	������{���B�w�������Ҽ�0�v��m�Œ�C�9���P�z]��c��?:7�$�i��X��;��p��ߪpHϻ��6E�g��,�����}I_ba�~Y��l6Q���-HqO�c��+rr��-�{ŧ���QѮ8-BE���ۆ�"�m��Y�����q�b���%��-�&˚zd�\�:|��.�jhJʽzi(o���F���g�I�(Y��8�r�:�N#Ӏ�cvV���*�\��w�M����,wƁ���*'�n9v[/Ꜩ�#��/x�����T�f�H�O���$�[�<EB�q��Ѹ��-�kKm|�&���.�3�f6p�K�k��̺��N<��1�[��~��ح��bk���p��kG���/���i����ro|.0�Y%N���Q��L����3s�,|���L��o0�$lB��o�f�}''�N׋,a|�8��_m���Ǐ<9��S�T�6��v�[�魽��#��m耛�����2��V��Z}�R���\�h���}��מJ��=*�[�4�M�Mǘ�
~I^��!���V�{�(*?ױ��}�-����s
DX5���ѯM𬧏�n|q³�:ٸ��b��h����F��+T����$�5���R����x����IG�|��ϺoJ�D��@x�����{%�^]�H������m�:�5��uE��%r$O�/�ş�3r>�e�*lt`�"�R]���L����#avŅ���}v�#?zN7�~gq5��?ZK]�Z�eI�͟Y6"7ny��1���k��,��Z��ц����Ә{��I"���=b�s�uN�>��X�ӵy�V���3��]�ӫ�[-3�(��,�S9���>�d�lt�7�SH�pR���s�q��h�#;G��P//��י%Sކ��n��uyċ�=o����������<aw�$��ۏ$��ƥ�����9Xw���ԁ�8y�^�ַ�x3���3����ݻ�&|G��#.N��w岀8��fI:��PEǭ}�rt����(���Gˢ7{?<���+1	h\2(���1K����q�{��������$aJ֚���q����Md�"VT|"w��5=��8����w�
g��yV#&^��m�m����ƾ!CN��]��y�e�x$��3��
u���}��e�#�a��[�	[ֲ�h�4bk�'��k��6Ф3+�*b8r�4����[�Os���Y�ғk������/�8ʩ���ۗ�0�I�@P��P3\:�{9P7�؄��u������I�&Ҷ���f(�`���<��:x�?����7B"�����]!�m��5�%������]/(\�x��K>F{Y�\����-�g�OMO��+�vm��^��nȉ�-SdA|t�߳�|}��y��k��C��B�cUv�;���\S8�v��{�^9x��
V�F[���;Z�S�΂ے-�J�]��:ͳd.^*�1W��(��xp>�q�A_�nKm��\�����k�L���x�m��X�p�	lm�Oɂ��r��7�n�<7�P��B���A���cZ��\���d]��@�vΦC�M��[���N�|W�3k�|���x�>��Ȗ�~���ܜ��+*�^�ؔ���'B��{U�s�y��	��(,�m���v��M�L�'�Ꝯ}��%v�ږ@̌��7(V���v�C���V�xyi��H��c��M��E�J��Oݵ�����oة_��7U滔,��\>����cA[��v�F���ي�C��t
ϳ�7�kv4R�x}_��|�D�S�Ʊ\�����8�5$�i�}¶�����{��N|lj���~�j �h���(#S���֑���\_#3�F�������я���dXN��U����'Uz�L��eq��mOS�}ۼ99R�!��SI�u���TkK�W/�w蟞n{�%�giO�b�I�Hī���5b�B���JI�,�D"ϰW�O����'~����]����4�Ϻ|�6�0�,k'^��x䄁s~3g9�0Ѩ��5)�w�g�ϵ߆T5��6f�����-~�,@9߳�¤��'�WV�S�1��$2pa�C���n\L��.�����7Rb���M��rE�n���TM�L��y?2���W���-.����>u�GR�G���٫�P��i���F�n�~�)�r+��f����O��/��ߔZ���Z�֢_���(a����s��w�R���2�f!q�Af7��N����~�ሸQZIKL�9��n���:����)���,��>��ǏÈok06�����|�ܕ����_jk_>� w1Ж��A~��\2���^�X��0�MKM�w�-�c�s]��{P"6^��y��n���O�5�oVz�&�)��#D��>I�7DL����M_f�r�b�>ب������g2x�i|t�a��ʗ���#׬Qb�
�%[�H�+�6d��i6�31^�:��"V�ÉꦻQ�����j}k�	I���>�Q��� ��c6��i��~WM�uY�$�m�Rn�運Gի�_�zn������Fh���r��Jϛ3�o����	�����V�6Z��ٕ#b����c�7�h���]��=N�ΐ�����PK�.ꤾ	����1F[��x��v>��2�oU����T��چ�C+R����D���ho��L�ot_����_tq�0_��qL:}!���G����?:�Ӎ�7�VP�=�6|��T�f��,@vfY(�hQ��u�<����u�lG��w���l�bc�k.���լR�ʷ��xã��^,*�� ���cO�i6~>���n��ǻ�OZv�})𰻴��N4(?�����'6�_l��J�"o�0Y��Nd=�'Ig?{�8ⓣ?�M|��^B��vٙ�� ��foM���)sU����	�ؼn,��.ʧ(Ca�ڒ��_(��%9C��Y]�¥�1S
<�1$�Q��6�mHH{��Dm1�_���� ϯ�W9�)v�gWT��㻪�n�	4�K|�:}<S;`J�r=�웒��e�[�1���ʱ��ļ#Y���E�����^����׊�_�S�m����I�8�1�Ζ7m��nb|�EK��mT�������Z�Y����:�V�=VPj��Z��	��Y(s��ܗ�T����'&��x�3��9�ۙ
�f�o��+n��f��5ii���oԖ�yc����m�����h�;�W�M�RSLD�O~͵�l�(����L�#gK)���,��NM���͞��^*]�i��u��V����%�p��r�=s���y��M0`��c���wlA�g�>:�"�~�>���-��bkl�c9j������"x����rk%���;�Y#҉74��5'c9�of�5��+WP���)/������/
(�8ѲuFu�㷡�I�S���U"kI������P�[k���v��%���뿟�	 ڪ��bf������� ��������}��j�r'+�l���C��ȮL�o۰UO\��kI��IG�^Ͽ�-�S�lV�a� �@nhCއ���VA�?�7Yn~�Al�����Y�B�"����R7+��ߜ�Jx��[��rq%���iT��'�>��������tۺ�9��}�u�wA�Ͻu�]��3"����>�L�p8?\{#�d���+�k3�
L�sCo�tX�	t��/�;�M�*��+�It�~�ů���)�))�:+�������.���^W�ǹ�O�˻0V6`�p*��O�6yi����1S�9ٻw���F�&�l�٩3�?������x1��	�zu�gA��Հ����}U��Z�'�Wj�I�b\�^9j�5&E;o�iK� �O�}7+Q�㪩�H�"W6�@����,���p�-j�܈���)mZѲ�n�͡h+�kJ�:�꞊Q'ҟ���wFS�LJ�ߕuq[���g�Fg��;�e9r~������)sr!���1���;1��p�����0ı<	N�8�w�ǚ/'�>g���jM2@��~,�MX����y��3Ѳѐ��������*�IE�In	�o���J��9�*��u�kO�'�w�HX��&�5�BdtfVůBl��^�ۚ"�^��ؽ���qY�����X�)S�w��`�m�ː)$ǉ$�\lo�i��� �x�(Od���[���}�8-��
=S�wEg�����pތ�b���G:(�+���q�B�žZm�� ���Z�$��&����\��a�>���X��I�8M�o&���H��?%��4�I���0�����=r��gwqd9 �i��ӏG�-l�!��]�À~�21��ө�����rh�A�׃�!bu���j���\g��: �J̱�������M��B�\�kί����XS�h��O{� {θ�����aMmk�o�Ų�K�Iu��& �� ��T)	� ���(UJ��EZ"%��B�P���z���<{����~w>��ɜ�u%�w���!wk�g��St,Qܕ���ו�jB^^�ڙ߬�sy[fg�Q �l��3��j�;R	TF3Ow���>�!2����0"v{==�}��CΜ_1���L�1�*pvmC�M��:v��/��	DE
9�� �����z��-�f��e�tA�\�D��kR�>��O^�c���v��'f �!�Z����X�a5٪_�pE�](5���y�G>���J��b���^�O!��	F���Z"�L�3�l4���-�c@�I8��y�S�g�9s�Q���l@�-<��b�?�a�؜[��y�0α�*/��D�9�Ȕ�Q�R|7��shl�`�����і�-��ǀQ����F9�KMֳ�;�jB����y?�����%�ѭ��'� �dFɂ�?��3�+�Kt����?�J��s������K��ٖũ��@��R�����~n�9}>�t�������{��^�'+!�;c�RW��\�|\F�n�k��FH�ƃ�跒�;Q�¹�%D/�jW_��N,�	�N��b?	0M�����s]����R+�X���gV��)�� �C��R�.�u�D�Z���7������>dw�'�/������<�׺��aږ��lap�ihf���L�nAq�@��֤�j� ş]C�w��J�#����E$ߠۂ��z �����|{��ǀ��^=s�Eѵ^ve�����C�`Qu�ÿ�9�u�}$�H�Z��S���7^�Y��A۩����\1���:/^4�%|�^���j|V�Ai��"�~����5���t\*���ǀ�O���9�������N���C���3�]��pL�=�O�[{�$�@߃�w�a��7z���/@7���5��T��ݮ�k��%lPgK���}IX��7NS�n7/�sq#��-�hN
@��X�Ԑw/W��<������D݈\����?��Y��l�s�B.�b1�G9�X}�°]v2PG�Ed���7[��	Y�V�74웟��ߋ��ܢ\S`��-�BL$ӝߵL����AkG1NU6�sY���F��%6�3�ԤV�Mo\N�*lxE��k`wY���B�9-�:5V��ҷO�S�t8�>��V��Y�}ZW����t������|�zL+�P����{��ZMdeL�Px-ka��`H���gDv�n����>������٬�X��$�M-1�Zߖ���aS�n���$��{��=|���t=���o�2�˩1�"l�6��"5z�uW^�lx�����63^�Tn����p}J��٢+]�5_	�a��ل��+�U��yv���xx9�w�
�(s���dE9'��n
H?2h�ۥFB��*Pz�c�>CCG-y�kt9Y�vm�@<���#N;ds�֭c���P���x���Ǫ�����d��C�&�G����d�����HM�Mb�=L�U��҈8�v����NGЀc,u3ukY���W��r ��!p�&fQ����p�G�:��Ф_��G����YGy�7���Z�+e^c1@��~�/_t4�v7k��`:��u���N&�7R�z�k��:�m�j��jD7������潌r�go��0-}��N }�<�T�����&���R^��e$V����|Юօ�]K�GM>~eO=ZJ�Q�.�<`U�3��MM����{���q��މ������-	N����jH����L����r���_�f��(}"�������8�4�y��l�D9��z o��jB)}tC�}H���"K�+�CD��7G2�lh�Wd"����{�����p��S��/��)�`G�sS�����L�+ON�;��>��y�>�������ث!��?�{5쥎2Z��z<��<*��(������۟�a�aHxh�\q�I\[E��9�w��slZ	�r����(�=����Hֵr(�z�ܱ���A�j��ǣ��0���8��[�a;��|�ד�V�$9ַ��U���R`���۞�n�qE�&g�T�I�U�l�&�����N�E	f�mM�[߭���[~�����E��^�r��u}I�5�X{���߻(���H�-��t��G��^_�.vS6dA�a���4���XR���:4?����>���#�G��aԺܴ���;�ed<�ü7���f���� ���{��3m��s;��qq�1ѡB�\�������\���^;�D,��XǓf�3��'�o=���]��	WX�C�J��x9��z��l�˴�Rj��x;��ԣ����v��~�<%�C�OB�|�Ŷ���g�|0�Ƅk
��s�1��P:'-��ϳ��f��v��\~��P����R�?.�Y����U��g8ɷ�U��Zd���_� f�"3�`tO�|�*�H`�n; *��.{�����N4����i̪ͪSKM����8R��߳�H���H��d<1Yl*�zh���[.�攖^@w"gaP�@f��,4Ym�W=�����v�g��_�<�·;�?Ģ�j�Ҳ��d��.��Oo�$���☍�ץ��*�p�\~���lQRK<1g+?��5���
����8*����Yg���v��D�W$nĆ0L#$_A��T�nn��`��v?�]�:��uv[�Hh��֭�X�iŦ̉� B>�!W��h�Ӝx��@��6�[O�HǀO���/ZvcJ�C� ���[��ߢ��Y8bK�5��F�a:"b[��8S����+���l
����"9٫u���$�,�?��G��3�תnǧ��e<�$����M�[�PQ�Fص�i��!K��o�V���Yȳ$�令�u?3P�6jd�����c��7��V�"b>&�eq���������lYJ����v>��k{&翖���hkOO+m��$=�.o}�N�)��)p)_��~�����%R�zԝz�,�rcV���u�^]r�]�']��Nq)�����E�	uO������]j�a�7#�q"׽��o��^�����8�{p;u�D�N2�eg�vl���=�&�2����ofٺ�K��%j�9n���ݨ��ʟ0�h=�̎Zn��gA+���0ڒR�0r�3�l�5��� ��~<_�2|�v᯸sJD�X9�Q��s��R��JH��HVp�5�_"F���hV�@0����w����|kʺ��uv�A�a}����p԰�^k���P��kd�*�D̣��O̽�8���lv�&��A�Bʡ]];[(W��hm���V������X�a	K�g�u^{�f�����Q�]L��z��Q��vFbh
�1��
��\�g@��!228bC����J2w�VE:+�[�;�"�e�if@����%jv��\0Dd��T(
,V�f��	�M��5�ƷV�n����k��f�d�c@4�HJ!����z�c֦�8ZU�޿~��j�y�q6��*��(������RQ{�(��=_����yOѤ�TN�U�O)@tS_9�ο������8ed]���f��t���6�~�Ly�E�4�)2�ʮ|$�h�"��O[���W�h���T�� �h����y�]�kNd��B>}Y�p2+3yu������}d��qH�D�Wvn#H�}13,D��+1��X������.��S*��\(އ��7�e�p�p�O=�.*v�g�{j��Zi�]\���6h�0�w�f\�4`�s/rjL����%q�?zҾ����8\ ��6����X�^���˶:I���3%�
2ٮ�?p���K��w���~��_ύV^��99q��D���{E��R����������?w��z��ӏ{��+?�����Ͽ�{��՛I�����.Vc��B*P���=,���8��s-3rH~�m�',���0?�l劷��J;s�r��;ʆ��������w_���!�.IEs5u�;�i��O��p��Â�����N�]R�O��Ub�R�'Ǌ倿�͵8�%[Oq^���l���Ruv.���wv�G͎s݆V$�8�:n�-�>i�
4X�$g�4�&�=�p�c�c�q���<uv���3�����"[i�8*�dSYG�J�$�;��hk�~���x2����祽rZW�r�Q��3�( ��|�/܍��Ͽ=E� ������O�����X����W�f����M_�Z�
o�#�B��,���
�������a�%B��	ڿ ������F�GAi���5����U]���Uzz֡��7-$�`�o���B@Pϓ�����!)���`m�m�@}�(�C>z^�Or3n�>C�Xm�۷��4L���(�^4�v�!����UwE-w���t'�:v�F&&��*�S)]Z�5�uT��y'�㺕ƻ��2�g����.g��N��;�*`��4��bk�����Rh�2�
�a���q/=N�8�}���K�?���I��#����|p~�������wĦ��0��(_�� ��+����}=_���M�BÃ{i/*u��'�B�����<�b�uU|�Y.�Z;5E�S7ަ�֊�E��n��`M��Iu+3d���O�#�u�#��:�9�F�tk��9���Ɉ�Ȉ]��d��٬˦���'��
7	���41�%�v�am!�}g������Ey-!�����E3�Ohm�c�r���o�4� �6����V�هG)�0�j��S���a,V9�Bp��z��v��}V]=ܧ޽��M�+f�K��;�[��뤺�jl�"��8�}gɉ��t�:�q�����k�Ź?�����u���n~���zW�ο��N<Cw}����=��%^6M���Tg~�܃S�����2�~'r�d�]�[sp��:����D,z_�g-�N�S%��LQ~쭘W�� ��0�o����YPi���{X"���o�!:���L*�~S���֜������7���xBQ�dxky�y jAz�UJ��@�	�l�2��^�4��������AR��t��2������|et�������@*J"Gn��7����?w�*���*���}��7�E�WM��ܜW��{��5�4쌢��HI�����R����\���x_�-s��<8��/H�@�����D��A�}��A�ì�*���v�Iϔ17��f��Id�&7K��*ͨg(�1od��J,�ZQ���g&���k< F*{{�+Iy++��G��Jr�e?�*eR)~��U>��p����٠9�Ë�.���ܺC�%����y�s(����Ur�y�S�mpB2�Z�� ?MM�B)(;�W�����L�����"�p�}��B^���vmBq�̛_�����N�B������z���v����`t2N�0��0�3�c�é\�ϴa�:��`�L�����Ku�f����
�7�OF��6�C&9�z����=�6�ч�u�WG���۾4�a��:K�?s᭎N�ΆGhIa�x���7m/�1E�5.�Ӎ��r�T���8�:����a��a1Ę��v��j�2	Ă�t��j[�A/>,y�ѷiJ�������>Tmj�fY����4r��������`�&�\Ap8��^s�m�׎Ӆ8�a�s��S���lU���q��L���1 �n�K��wSweҤ}A�.q�n�,���������yxh�6Sb��I�=α�#�.8{]�Y�^R	'[V�¥P�5b����{h�T�K���j
��|��o�	��6l(���U1,ߋK<����g7�M�d~���Ϳ���U
1�H爅p� ��9C��^C��SC!zi�j��fi��	�%� U�d�\�MH
���g��c�Oc2�����b�Z�N���?�6�`�!��O���;`E5������S�|du����g�T��3,k�c�����Ǣ��N&���2���Wn�󞲶΀�gH�S�"�q�o�(�Gag�I �J2�����  ���י[cR�ӐO�ն�^
�����oS���6� H�&\�m/�b17���D�Ϝ�2X<�@R.�	���q�\,��ı6T&�Z�	b<]N���$��LTHs�%�U��Ã��Gsyc��k�Q�P	˝�oKs�/�m@�r#	�����l���*)��=��e������rF����=n B��Ԅ�����d���(؅�y����J��2}���>ڣ|q�R�ޚ9��*4%��sC�����;�p�������;;,�a��p�Q$�����>'��;��kW�S0s�"�	����b�̅4����Y���H��o6�[�G'Ze����n�r�
�2�� _!=Рr}�������H�X�&�N�Z`�~���[��K4�f�,ۣ��G�B��]�&*����N�^�Q�3�B�v����v�wJ�]!�~~0FOI��e����6�犔���%�5�ah��N�1`{ϝ�,�sv��
]���� �<;�u)�������8#g�~�9����q��Oa�����G�W��Hg���)Q�d �~������N��8א1�Ӊ�:�>��3�!�ɵ�}ȧ�a[�b�8�gΜ!�=A���(�v�����_�΍5|<�3#�\����]gj�ak�tc$��z��"��-���,, R��3�Zާ���_H��NI�~E���.�#�4/%y�>�t�e���˦��G��
xi{�Lq>�xT��~�|;\Ew:;�H#�<8��0��ɾ�cW��l!��3�zx�E14�d�:����=v8R�|e�GJ!���`�(�/���2�_�p���g`�L�����,Pc��A9�u״瘿�,��t�GGgW���5�!�0�v(;��FSq5�uBiX��J���
�ݶ�~���?��5u�dD��Nh�w�kEU��HB�E�惬�ua�����#�r���YW�5vlQ;.�i��oby>�q?3���J*�B�Jv-0_|�yd��_��,�����HZ2r�ѐ6*���;�6�\!o�z�,��{���#�i��:C��ME��Y��>���we�y:JŅմ�;4�ތC�,*�m2�7�þ�+Moװ�F���0���A��]}I�/o���ѝg��@��O�O�9�<8�li=벻BG{F%� �mu���~��5�>�mp�6]��&G���{Y��&������
�V�ǀ���U3�2�P���H9��<O'��	Q��=�|k�QuB��NÖw-���3�?��!�NTp|wVo˶ה��~�d1�H/RB�F��>x�}P��O��r�`��O-�h�11UPBOl|C����,ۇK�܇cӿhj�g�q�ڄ����#����Xi�1���f�Y��.x]��"����:1{�� z��槓9�GH�ڔ�5��zo�b�ٴaS⇶DL��㎣�lR|�d���C9�_�da��OG;�����$��V�`<ȋ�k�_��g
����!4ʹU���d	v�ggV�����i�?Yu�o�3�Y��	k���l�ħ��������q �Q��X�K,p܋2I%�l��.�D�i��|m\�v�lΗ��*&a�h�DdE�$���:|�:�`��!�quݸ?0dd�50��\<H���oM�rK�j�Z�R#%<R�Q|���F��x�N�yD��}-���:O�)r�3e�)�$l\�j���{����h��=L�<e�A�G���f]������B���zZ}Y�&�pk±���5C%���)�9�\�Եv�0��vIg��'O�xl��k{�l�^�C	O��0��b��系��%G��9�������u�m�^_Z��3�:���g(���t�x�U���jx>^�:ϩD��K:���/@��}[�s���(gȝ��GUy���^
�7�W!��t�^q��I��E{����Ժk�m3e��#�9g���r��oh$,�����t��n��:_c
�(�j��*��S%��Z�Ժ�
-;�kM!4�#��F,�a���˪�1�6e�㨩[�LV��d2b�B
dxf� )罐��63�Jש�e(6m����_�}�>� ��<�����&k!7��'�v�آ���?��NR1��gj_��t����7�@`�ta ���cgnk�*�������E�]��}Y�)����1��0|	���5I��6C�fos喤�2W��k^;�c|o-i��S��[?n�ފ6m�K�H*�/X�H�l�n4�z��z�]�>�P7���|��ݬ��-�p�[3�N&?��3��C��O@d�نS�b�����J���)hb-� �0|o� �9��n-�P�d����Y��6-Si�U.�dt�:6��jV߸��|&	��%�Cug�$��������5�;��F쵠�0u�5!O�����������tg[����j��������9�p8�8 �����H1���F�S���F�|!ʥ���M�Ϧ�5ICe�0�`��u�{1�|��B��P��B�W�o�6F�q!����m�ֱ1'C�6��/ݧ/O%�tN��g]ڟO��Ɵ�lR={��g���+d�2O��:WF^�֤�8�u�}���L9(� ���4�_T�_����1A�����%s�yP�+�m�D�f��xU���$'����_#0���ɤ���	!��`q�}��
>[	Ϭl���v�!5���<8�dTD������@��gxx�*�h�)��f6�I+6��7�H$I�߿��4~U"A����WM�ߊ��T<�{(�����[mcj���$�c���<j79�(�nh�������KB��T��5� ���M]<�C!σ���D�w�Lr�f��y�ݗpq�0��k�RU���>�9Խ�xX��"6���q%b{��ۭ�}����B!iq#o7uа�`e�,�+���H��=��|ݤ܈8�=t��;��A�6��w�`��F������J�1�����D`ӆ�
���{�W��<A���!�G�0J���J�
4��b��kinh��T؂ [��i�x���K�>����-�K��j�/;	0'������(˙�yu��1/˻K.P-|)�?,4ڂW���0O��m�H�Q����ͭ� �\,k�;tZf����'�B;�'�Y��M�Q�cXL*nEء��8Ad��%$۶d��s�P{����\kU��#�B�kK�eEx���7E�Q7���K�Y�6�l�����v���"��N��XJ��:�o����G��D�I��j����k_����t� �?�$:wN,��Y.@{��N)0�H���4��3]�8��N�a���J������}�h��a�|�^�Мˁ��íi�OiV&{_ �|{�$���	%-��>ƾ�ϩ�3���s����kN1g�|����1���ڤa���!��v �|�C:�"��t�b/�]�;+X���K����=���*A���	�DT\��C��7�n�$�ٺ�֐Ѝ(A��mc�qvп�����k�@4֏�&��	2z��zd;���^s�U�ؾ�c��N�8w#��ܧ���5u�P�������'}vj�.�+_^7�d���z[G��{���>l�q��� ?{L��_7~ˆh_��
>i{����&�.���&���,�77���Z��p	/U���ę��R��vI���� 
�$uq��Zw�,�[P��Rߩ�})qi�HQ�*0�@���H&�<���-���Z1)_�0���P�"D��9|�vP�i�OD��P��6�5��e:�oZ6LK˦�Q�fB�1���)��q�6�Z'��]V8��N�)A�n�Ď���~eN�����B�v�6ի�w���[��T�*���R�\��I^ouPwظ���:�>~I����@ZV�*�'D_�A4a@�d�D�f-�X,��ˡ�
No�&k����5j��`���#h�iy�i�[祽���=�=+���yj.�d�8hY�z���{���/��'�%����B�?u��x���=FU��9�� О�)?�|��l���X�B�:��p����
O���Y�	Q#�z{�|�1�j��f��3ck��<j�KY(�K1W�U�U��B�W\P��n���b{g��PC �=y�I.�4s�ο���ݐ�&����?*��"2�4������4h�����`�������&�ny1o��?g��j���;�@X��/��?�Ӭg��4)ɦ���R��In�?>t�e��E��,6�.�~wM������$Oه��8MyE���c��x�!SZf���\hI���Z��l@�c��:  �ϫeE5?;��n|n$����nǁ
��3q1�����
[{8���S/ѣl�h��N[VԦ��k�!�;�Г��E`���e�W!����9�dT>������p$�<��ۈz.><���g��P߁!�����<J�&����Q>�Y��Uf��@��a�B���X��x��T���Ro�W-�ρ����F�m�,�$Hq���dr�K��̤�8)�\�ɯ��P����i1ق�ֵ)%�z'�������@�;�_R���h��;sґ6'/���$���E�eyu�vN�BDj�E"��l���qH�cF�鈜�nc���͊/�2�E
;�_Wŗ�4���9Q�ki���g�Cv���s!�5<�#FJ�QCSor����K�P?dC�S��y�;7\�W+ـ��Wx��:��'�Ʃ��巶��N��Nu^���+�K��gF�Mo ����O�3�RMט�N��y�1�*���_Rvވ����*��r�x��]�1���t�*/�ܫ� u�F���1���`<:@7a¼�Y��-��|j���h�Y���y�ZH��7�ڜ|KЋj�k�{nݐ�hSW���5=wb#q>����$>��DG킽ݨu�nnu�,��'��^���-2��CJ��)��r���(��x+Cs,wV�h�N�ƨҐ�ܴbO�6u��u�&��2Rf�����Q��6��8=�k��B݉���z�Ѱ�b�R#�r?n%"6ޖH�}�LLx��{g�÷z��%�s��WcN-�c��l�D��3e�:8�4<g�+�;/�k��9�������1]-X]]Ȳ t���)�|$���zgو��E:]�1OW��`��+����ap�y1{�m�eF�M�x=�����WW���G·¢+��j��oa|�!�����J^��Ӳ�+/��4%9��54'JΚ��ɷ=KJ�H0�/�j�Ƹ/�r��|�_�>�����{�Gt6Nks��H����Yd/�޺�k�,�A,��vK��x�u�(��Zd�8V��a���C�WN-���C��L3�_���ҝֹ4ح�&Nl����v�=j=��ٷ�M��n��(4{W�t���I�v��kQ6M��
������
��������S>Ua>���\���W.��~��WO�v^�3�s�^��u:�P��4�r!Uy�_��ZGD᧥��Q�Ł-ɦ�e)O)��Fxԕ{��h��I���Go�Z��5�����T���ϭ��%JK�:C.���Ԇ�Zz�#�_]�������N!`3�5�%E�%R�W�@fX�aw��. �#�	�7�� 3�u���~��t*W;�+��&���<��;�V��eS�Ʉ�P;�`�+��~K8�=*h�	�6u3D;u���x�ʷ�K��d)�Y1N�D.�M����������1@3�<�]]/ê2_bp�&z�[��Q!dn�Қ]��YN�⎛%u��F��Ķ��y�B+k+c��Psd��1����L1�~�$o�DA��D�<���3�ּ������K�3��{!,]T��Y�͑J���'<�������l�)/���׏F�ǀ��f��Zk�aY�A"i��$=�v�� �Ü�T�ק�߻ �䲪���ϱ��r��(�z�la���g�w
������"b�g�������f`���U^��c�\o�X� .���L�;2ʢ���D��ai<�}y�ک����e=*����l�c�~	��c�㹑����5�n������A���],��� ޔ�QV?F�'�ׅ�Sor��
��b����aj�
w��܀�9Ve�-v'/�-H	�q���ru��ka����q^����vN0��N�y�iO%�u
�� ��,��<>�ɤ:� �J��\n����1�O��ª�����&Z��&��B�g��z��Q�H^������B����V3� ����΍V�iލ%�t�$�� �4C5� �4�D�"��I����DR�s��W5�Z�K�tE".CL�7p��(��=
���^!ԡ��'��"Z�ϓ����)F�K[=v>���/k.�G$�<�u�S���#y7�e�$�#[��c���1@�P��`f�n���������3KQ��m_�+z��$�)�$��̓��c�EK�C�t�V������!�%���9t�E̮9��Ͼ;ؘ�п���n/R�i�}:�Ia�1�+��e��n�Ű��C]*+�WH�+M��~Y_R�����G	��Wyh���2E��T�ι�/�0�0�Q�3�����1C[R�n#��DW�4���;6��n�s�������AOex)�(��u͘D��c{H�Ƈ���~��lF���R�U3r�������Gzo����j�X+M�nY��>��f���F?�G���f��0EP(7�ʳ���{�,�X�����q񮵨�[���p^��Еi8��-ܗth�^s���lk�z3|WRu���[K%ݳ��8Q�+���"�q�U
�Qχ_���w���}:�T�J��}P;� ���1���s���Q_��?��a���gt�����a�]�X��6h��J�S���&��Rש��i��m��^Z����g��'�s1'��s��z��d�t��X�H��������.� ��Ij<���5E2�Ozp���XLW.]��1�S�h�n.mJd�O�L�H�n�>���!���*��Z\�he,�Ĉ0�b�m$Dz:�Hw��I�W�Ki���� K3)���e�eJ>Q�iz�o��1��71Z�#�r�yD�AO�򨠶V�m\L�X��*��s�r� ��C�5�m9�#��R㛑��T�	剒,�`ۮ�����ݔ�"�{Ū��CV���{QƜx��`��VpC�~��E�, �����}�C?�q�W�Vj�Ҝ*֚��-os��!�bh���}2(>�-u�N�)���9�y�0JQ�0���gs��$W�{,�R�->ڴ���+�iYw��M�L�ƐtKl5��<ҹ��H��q�����	?�.R~{
ѧ���Q��q#)kw��f#�M��vsm^D�hhmF����5���
�
�OX�۵��R�z�2�B%�*L	�)�'6��)����}3]L6�ut2MEQj6S[�-�V�2P:���\�D�%��X��6L�z���Q��t	���T�6���Եgʐ�ծ~�=թ�,Y}��	{�%F��a����`�����
xP������ڑŽ��u����X�AXi�f86ԅn�Nڼ�}c~�.QE����2^�n:mࠞ���sV;Ӏ�{��W���ݙp��O��J�g�,���1���Ic  �' �'�>��:�زj@����B'Q��e�7�������������)�!�[&_���zH��(e�R�(���eij~g�Ũ�4ށ�y{����oѻ�{tM����"u��M�|^�b@�7��UP�U�k�FVX��T��W؄8�%��hcB��w��[��̋����޹�x� �6V�֞Atß������z�b���Y߉�8,�miz9�h!�冭�-}��U���/�.�r��3��%��
�f lq�-��ި;^��.i%*����1ik?�_[��t7�*Z����[;:��tۅU�L�b��+���^�l�#�	�_�ր��F��|э�\��A< k�!�#veI<?��5����s��ష�`S�q[��F*6��N"��uJ���|wذ�[rT�\��&��O�^&�m���$�����q+����E��*k���8�P�U������1N���Xe��luw
�f��AU��S�"�a�����l�GI� �Q���BV�˲���m�T��"E��ӈ�8��ZqZs"^������B�\:�P��=�gǗ�@x=,��ٯ_Y�'H��Ɗ�?D��F�J*���5#4G.����gD�a�L�M�X�p_�#��@ݴ5�Gk�l
������.co��G����镖9T�V�r��Xa���Y���PR��V�a;S ��:�u?U~�{}��g�/�=�E��
{��뗣;�?) ����-�HbYY��K���j7������h3��I�D�utA��נּG��kRŪ�q��%~�hzB��HSOq^�jO��"D�Tre�Dv�������g1z]<���V�璐k��d4�+����(��l���U)ۥ��'̅��-��������Yx�vFIj,�A��@Od���>E4���\��|��f���ܜ����M���j�ń�ѯl�E�1>�_#���R�-�8fӯ�HK�BT?͑4.�X�����;�4�-b�4T��2��z�}d�h1oĞ2�?��vQ~�~]C�a����A�X3��	2�ʂS�f�����	%�w�؝�MW����0���޻'�K �F��cn�@�DZ#G�*����hc�����Q|�!���B��@������M��wSiD�k7��IR��M��y	�X<%ܦ̞���A���f��ox�o��4�jB��0.6+����dN	���l\�I�"�q�rߞ��
v�Z����ۃr������˄����4�\��/�㹸�Ap���fM$~:��_QF�uCt`#�H�+�gn�K'�;u��Ұ�|���7H�|"�WOD�JӠV�b��8c{�-q�X���)�k�W�[z9ς�!�饊��Fؠ�	1�q���N�9�j^�ISh/TߑJ�
�e3sa���H
��A���?p\�Xt���t�xJ��b��"��K]��7/����:U�\��?�6x�o���.܉�|��k�̣�C����K�~����Pp���u��6d�;�m�HQH��4�*�q�)6�/	��*I�H������wV^d�r���8b1�B�h�cy��t��6X�i�T'2�0�)1��]�	� ���X9).p'�;5kK�Sجm�'&(�R����CS޹��Hԭ�T��ټ=����Iע��8�V��:^~5.~,��eC���6�js��Jp~+��
�1��k\.r-�]/�2RZ�'i����ّռ�h�����K8\�E�~�Y���]�|���V4��X�kR�W�Ƈ�����L�Q��j�R
˸�"S���ޝH�e�F�6`�h2O�Uz��h��$�˘ws3�p�% ���b�b!X�N$	��mB$�z��w�;�į��# �����@�T����üP"3e!��e ���NM����d�e�'���u�ru*�~S��e%�����%��һ���I�A*�z�f�J����8z��fFO�d�`UM�HJu�z�RK-���HC:h!Q�	E���fzr�4���y7%"��C5%�І�DS0qy<���H߈.�Ֆ�u��1kёО��������G�0w}mHd*�t�Ey������5j]����*�-�31٩d�g�����m����"��D�u.��""�W�|������&�P�]��#����z�<��X�)�Z$&nK�mq��JVX�̍�|��eZե��N�=��a��(I�K���* hw�}�ˑϳ.x�Q��r*|������\:�����'�o�`31�ɤ<�9��Jq�|�y�K���{�
������/��/<%GR���Ɨ���Ykb8�����"�L)p�"a���:�
ΐ��<`�cր���:��K����Trx�z^>�P�z����: 2��8��ꨕ=�N������]��C�Ïy�����-��HgpE|@������e�V�V�-=	A�d�����Ԋ8��,��O�O�tvŀ,Z���$���k�P)O�j�y��q�	��xp1CX���"쌲2�̊��nW&L&%,�ρz��-���7%�1�v� sw��}��h/��J�rXo�t��s ��QA��W����:�^�=gXu�hW��T+��_��u�u+l�۫X`�$z$��@Z0)Ʉ!�ߥ�㍟^��x�1ksg�i��������������
u��C�Ul;����&���1��i���P�O����%&�z-eQ��먢f�|����z��&��v`�ڰ�-��E=�`?�wǀ�R)F�*��|_oD�<2L-��CUn4�f�����`�icS�Rp�L�Ƨ*H�� %AP`�-�̮�`��6u�zM�0���z�$�;���
�H�+�H��t��������'�.y-:^�u<ˤ�_g��ptj�����JoMʬ_�e(�U��P�wkx{F�L�؞�hɼ�T�E���Tu��,˾��뛿i�)C3\�o�Vq�5M��&A+���Ϻb�S𞗎V�`~�%����g��G���w�3NG�} ���rd�~?����;�J���L��Ĕ�1.8xԻ�ms\hdxj�϶BM�d2"HϞ)�2��%%#� �M7k��6I���x�-�E��Ue}y���b�vZ��517C����X�[z�O���bȗ�m�ݶF&������0s�'0�F�Xk�G�Dߌ6{�/��+�4�v�F)'{Vy��ʊ�$#��I�[�L��wI_���[݅�k������=G�m�����J+6](�ڛS��� 6�j׈ Fk1j$1�*J��Aj��Ml7=���}��ﾯ����#�w��������|=��+��VQBh�{�⌙n�^Yz��3uz}��U֠N���H}p��J"2�r�J��.+e�tn�X�_:d&�\��v���m���K��`���ik2�37�M�s1���Gq���KPb��y۶��\�B���s۳��s(�Qu�нj��8�LÆ��ﾰ=+�L����s6�Ϝ��2�@��}f����JUk]�?�m���U��5�lb%�}�а���j�U����1=5�&W���˥�t^��!��:�J���<��y���^'�+��w���Z렘�ʫO��O���+_K��wC.�J��F#OiKFJ�+�K��l-��|�kq�_Ķ�S7�����̽�#�Y#�i{��
�Իn��cӔL�R������=X�j�ݟ����-]Ud�4�є�J�=n���`�����]4G��j`��v���/0��d�����5�H�XK���5�S9%K"�{L��؆7��g�$��E�l���WG\��Cޏ�#|���_�)ǧ�33	��z����r���B�{S��?���;@�Hԛ��$5�ѷ��9v�>(Л��^��+c���M���)j���؆��.��Y��rU�[� ��ir��]ze�䟔���KƐ JEP`��k�������}������!| 3=q8�.�w��%��\@n�94}�l��(�`��ްKN�N�9��L˹j�6�*3Fͷo��\h_����IN!�O���\zɌ�q���T�W��b���Em��.�8dp��dI��k�]�]I����C������\	�(݃�G� ����ے�ՙr���Wɉ��i�m����=�'���ĺTH�:#�)�h[�G�Ф�*ׄ)� r�Ʊ/�cᥲ��۷�,Uػ.��Q�D6{0t������}&ؠ��2`��В�m( �yN�f�J>E˴i�i�/f�{Rw#�hS/�ֵ/�ze'u�
56맴��*�/���ϻWhG��,�Ms� 𘚖�X�;�Ui/Y�O�s�.���S�����Wʭ���Ǜ�`�YD���rrIu+��*�ܚ�f�Gy�����ehF�`�T;?�)���՟''��ą����,G��Y��^��Dw�J�X@�˕��:R�W�{ҥ��&0����^�371�Bsg`�`x��w� HrS*ަg�{w�V�X�Y�R�Bt�E��Ӊ�����`e5=��
%�E���恧d����8\:JDG��G�c�&��c���;Q�/l�t���p@����@��l�D�4 ��m����!��Dhy�q#������8��<�@�pIݤ�5�7n�8���f�{�sh���[����F��;UyN��:7�Ӷ�z�ki[��� �9�w4�x��\���h�����F�E���vӠ��`�#|b�:_7��]�2���B5F���^�S��O}7�ձ�.OȲ�$9Չ�`��:JS�I"�V�Rﶲ��˾�E����A�����I��B_'H��Ix���u)l"Q�E�.��lەr�6ګ��b=�x`�^�cQ��$jW��=���_���K0�!Ę�5v����_���-��qױH��(��n=�)�kZ�����fŞ�儯H&���f�8�k��7�
��+K��-�5w��mZ:�9E����0��vE/��n���=|�{IRi+q�ai�qu�,��75��L^��V��v3O�Dy�T�|Mt�!���	*K�1�NY��оg&Ȧ���'�����l��F����fC���ܴ��=��#��II���r�M�O6ꔔ�KZx����{a�/c?���8����d�4�-�dg؀�
�{�t_�y�8��-k��hc��^��~-���Ȩ#����cӟ$����N.ڦO�C�Q�~���͌^�.����w����h�V\��b�F����KϬ�&�u��������z����5�'SX�~l�ز>>cb?"q��i�Ƨg�jO_��?�ǾY�k�~ѻg��iS=c{i�k���_��N��X��ν���X	v���3���:X�N����;O*��?�S�2�KIHK Y~���l�}ѱ����@�r-2���m��!�c�_\�S� �n};n����ө���{؏���3a@-&yH�t7��y�Sϧ*�;�t�u���\�4�@4ﴫ�k�i2�߯,�n�^�H�[�nk�����K��;�hC��m���7�������w��y*�}k:��W�c�^e��U}�*�+�A�I��Fcs�-����l���3�q3I����6�d�xj���ui����.�ת������"�6�ZQ{�*tF?`��;+�ႂ��,}�'(�_ڞ�$���z	�Yz��yC��_B���RZ�OY���[��['��b����?C,�c/�V�YE�^�;e�ߌ���0�j�e�+��^���G��M]��	āG-g�y����z���Hu�1�dwٴ�Q���LV)n�w��fW㵱xĊFEf��G'.p��n�h�ܗ.����]�%�X�4�V�k�B�3�~*�~���&	�U/c��o��;_Y=?�H8@�ͤ��^,
=*[����39��Z���"³DG�kP��Ii����҂����c\!�@*w��o���b��_���C�R��ed��Ns��O�A[h�/_R��R@����~T�W��*����)�������G�N_3�^������h�_��o� ̀����k�؄~�6;��ϯGұ�ha=�����q.�w0	<oU�@)mj-�6;H
�LE�_pt>�8��o�nʼ�֩'x�7��|`�r_�)�R�%+��3\pr���3�mX����RJ	�>�xA��&,~������%��Z��l�8��q&��ug1g�H�S_�fW������F`�j�m�%2̍`�@|�5U�'�nKCz�:,vt��)��\��hz�%D{*u�~��g`�o]�<���wJ� �֠�����3��Ô���R7�sL�I����3����։\��ܖ�L��k�_gF"xrh�m��������d��ӅÜݶ����)������_5{�
�]��2�4*�����}�%�� �#���sa��X���I?M�xJs�l�X3Ǎ6n�������P����Q��!��B��DӒ�t��~{�Ӈ%w�~�ev�N�U���\��έ��QB?i������C����}�ԇ�Xu�$�V�A]�h7+t9!��$#�x�Uۇ �dqF�'�泫b(w���!ł	�3�		��oAB��q�^��*�8�����[Uy��ↁs>���T�b��{\�uG�
Q���>>������O�����;�$��`$�Un�
dٴ(�����x�i889z�.�f�C9�� ���j$�I>o���[F �">��N|&̤����I-�`,>�Q1�)��^�z����_�� �����?�\������8�C�\5=��P~����`�h�p9*&� 	5�� E#�E�o�;�v�h��Y�%����SJ�&w�F`$��E8Zc/�%��L!k��ln�"'��<� �QH_��h��z�ʈ�ݕ��8ܾ_<�GN��p5>��'�`_�	��L��*R;�h�X�~!���ڟk������gڬ䃀d7�K渡c���,;�P?��!���Uq{�j;\*��zw�1���߱Ƣ�:A��ɩ��}�DcZ|d��(�U����>���u�ْ�_sGϐ���maJKΒ��4�e�MY�7��W�F;;���oY��8�5[�B7
�^��_�7���%� �o��ub��>y�m��|�04T�FJ�R0u!���Y5�z�����xg�p�M�1�S�Eۥ�/fϪ�����m��~t�LB�4Ƨ��r���
���k�쀥wN�9׳���s���k\Es�H�Q��K�q�_l�3���#�N���n�~/֡��z��'m�Am@��|g1�nO��_�a�E8a7����!5����&�W՛[�A�m�.>xôO�)d@���&�����G�w�����i1(!���Vg�WL�c�i��gX��m[�/9�n����;��m��tT������`�
d��{��	I2���)Z�Έ ˡ;�J!gVKaԖ�l7�����<B��'�Z��7F��O�e��bm�BƏ٘��(���7�� F��n�ln>��d:V�oU^dQ=�;��8�s�{��}�b��Ž}�~q�(�na����� �Աb]S9V�*�'x���B�m�3�Q���ˬDh]�2�>:\;l��9@A��/�|��IQ�S/)���r����ǵ��	�-}���m�d`�LzV�$I?x��նb}�2b��l2�����5���k�RgXKZ�g�?��r��L���.��S�\	�f����ZM��$yJ�Z�8F���q��](�1J�ݐ�o��W�Y�A�:�
��_Sy>�Θ(�����{�o�K��a	�Փ���W[g�EU=�
��y��	$���ߔʢ#Y@��q�9��=,x6�1�P�B��j:�8�!K"t/!X��׊��@��(t
Pm�{��h�Cҷ�vN�~�,/�zn�I��(v�
j���l���l2�ķ�#��u��� ����|��d)�Q�#�f��X8`�}�Q��@mD~�5=��T�v���C g��dϜK�TG���� ����f�Wj6�-��Y�k!�CZ��u��j�¸$\l˓��>i]�.��H?0�iS�������6?�@0(T�9����^�l��l�-��"̕�zF����D�����ӡ���|��g������բ\����@�`	\��p-;�鶹���v��Qs����ۇ����Q�_���7l�/�Nf���|��q��(3�&f��g�݈追����U��`�pT��mok�t�&��\40�WPm.�m`	�ھc㑙O���0������B�nᬮm���w���JNn�8美�J'	>�K�1>��qrzW�N"�H��\��ͱfp�F/���3��D�N	�e���o�M�[�d^6��N��Z�_�tΔd�)|��k���bbh*��lS��oԂ�W��z�շ�]7ѵ�������G��T��P/wL^j_�B}gȻަ;��L�}�~�{k(-Y����7�F�^JnɃw�t��c���U�h��+����D�����#�q�������'�.x{��?h:O��mC_�1�y�OAq���>���ț�1�iN�i��>w���[�
ehO��N�Yc����2�}4�䗴$$�iJ#�zӮw+��;���-fP3� �ٝ1QT����dYqZP7U?��l��o�E.n�kӡ�P#ضX�W�N�>Bن��p��,���G�,-�b�Y�O7��cg�Ĳ��%��%���VF���KE�"g?߫*ŉ��Vɨ����)u������^Z�%+��*9���؍���ü�/K�����q8D�a��E�ޣ�9k3ELm�\�z��U�iU��u��>�74+Ϲc�w(j]#��Ԝ�����'���>�朌`:������:��&����E��ݱ�	������g&~?�٧��c_r����S:81�,=��-��rE�158�^��x�_̊�H�aC^o�m�xd������8,%��3T�N[mŔ^������[	v�岢����ϩ!���޴{��ԆL����7���Y�i�
��N��[���+Y����/_vk������"Av2��:�6�K�n⊌n"vT���v E>�d�j,��	&�g0,[s�<@v���.Ŷ�'�����Q��FAV-�����.>(h�Ƕ'�8Χ�һ�J&�1�4Je��V[�����=������n��Ξ
A��E-�ii&�n��i�Y�C@����I��.�[ta炄��#I���s4/����ӫ�8ꬃ��}�R}g�fZ��.����p�^���H���*��=ەz���j-,�����D���@����z�p���ŤdZP�Pa�xٝT�^�\(��*@σ8$�SY�KB��x��A8i��N�B�[�����e��f�]����2']ۘ��e�Ûu`jȣ�U\�?�Eӻz�L��`M`�+���lK���y��?M���m��W�����%�:�L�5�K*���{c��F�Wg��x�UV�Bo3��j�a��V�9�zg0�KF.N�7O���k+՘<�T��ɞ���Z:u67RP���='m�p�|��IQ6��uQ칐2<-�<:ʒ���Dj,��&�_��O<�:"�R���3!B ��{LC�V��m!t�qb��A?l�ǭ����h�4��6�OLO��;���	-������ڵ � '_0g���]�O���'�����6�ơ�5������
4��f�{�u����lh�P �[$���b��hr��ƻ�ˑ$�g�(����#���o�u���X����Sc�^�=Z�)9���i���7��Pꂅp(��rtފFםt�Z^��
�Hd��=�W���k��(km�@�	�+3�e�FO����j{|���4��KZ(t�6?:�O-v���sbr!Sir[�Q�=?��;�*�n��b�"��J�7�f�n�$^��R!�۬Ze��Q�g^�أ�W�<��f�03��x���8b�%���ݼ��]����9G8���@�*�;1�A�ot����"4�F3S�[B@y�%]�ۭ�klk˝'j�|��!flYi6�����|��^-by�z6������TF���Y�!@ɯݍ)�T�ݳw��D����X�ՑCA4�}�).�"?����
y��K�3T�Y�wXQ0���.�x��a�&�u4�h�Cr��;��Qn�C�����I؞e�b0�V*�l�-y�|:���4��q��e'K| e*�7��J]T,^Hϔ��,�N��=�L!�;�&N#d��[���._f��+dj���r3zF�k��f���S�%�m��!����zJ�R�F^'(Uej��*�G��N�0�2^�S��Cěс4	e{�]UN�Z��i���x��;)_>:io7�t�3ADɋJ�B���9��x>Q����&�݋p�C�P��2_��ht�5,��Zf��Z�O
��N��`;*�D�8;��Ε�A�� �H�Px�$���ܳ�,b���	�����䯿�/لTN!��"����@��k=C���5?�h�;�>ſKSF�s@yːL�MY8�j5��S�T���w�8!5��%�#/_�㎶ؐ�Ԗ5&d����ݔ��tc�:!QN�fŬ����A�+�ɷ)r��p+GvL�nM��c#�(�=�|8����O)J��Ese~f���>�[�E#w8Cq��c�"�"�[���%y���.���Vr�_��|�Jv7� W=���s�O�}�ɺ6��6��R;��b���C�XT�IP�Y�� '���{&�;'k��=+'>ʛd<�bL��Ib���G�P�́�IpZ�ӈ�����I��K�aM�o�Z�ʐ�	�vd���}�R��|� ���<���-G�e�xSO|>
#��1�����+WL�S�xj��<8���s�?�an��te��*�;Ԩʗ���S�6�?��*d�+�1�R�c\�2H\��z>=1����ad�!G`���3�s��P���z��\���\�}˷7Z%���=�tm���K�#���փK}�ƞ"G�3��3:��o��o`;gpB?����%O�NF<�����ڝ��n�<�S 󥝣��oe��_��qq<�cۥ~(yW{p��,�����2�,�:Uu :�~<H�^����|�l� ���F�%��]%�T|K�E�s�/ɴ凗�h-�܇�enT;i��-{��*%D��7s�ٹb�!��W���tꚩ}<dqO�J'9{w��͂v�Y����=.� ��:yW2�T�]gA�?�e���!�C1�&�mN�\��ɫ~��Q�`	���i�^,�,��%O=+�b��$��:�t��;=��X������������.��j!l�>�����
�c��a�]	�iJ�k��(�
ˠ���ZYk3��ZeO�p���X^�L��KtT���k~q�A���=��������ޮu����P��v�Bl�M2B	̝���ؼ>Z�i5�C��@��Qx�	�/j��c4S�� �Щ{0ʟY���K�T��������S����:V4 ����U&����\��}��^֒M\���v����$��5�%c�"��zI�{�S˲V�kс|�#�����D��d]!�'�G�&�N�ɡō8��X�/]�k317f�H�DE�����q�p�h�t#W��/34}��/O��j�}q�[3��B����0k�����<c��v�|0a�L/]qgS_QF9S7�u�=�v!!�$��Z:0��_������+wbl��*f�
r���.��T�~8����EC<�E}zO�H�+ 7�y!�Y�.;|���*���}`���W�=��VL���{WM]	�Z�C�0�xf�obf�{�%���*`���!@���	u�t.�i����Ւ��C4Q�`��H鱏���X�ch��/�����b��<�-�fU�HD�JCRso��9s�)�Z{i�-��v��]�޽^���
�}�K�a]!�y{��Q�N���"יBn���a�8(H�!vr�w�7�G��Kx���d`�K���OI^��;)�(�n��2<9���m��+ٛ>�5��2 ^�Tv��yh#��_ъO��F��[.�/��!`�k�Iݑ}�i�0��΢Uᔄ:u��;���炊Y�;��W'�'rW���%��ɤ�@�Q����!�;����g3�B��T>�4����(�U�&�\
n
ba&�,���e�{_T�#s��4�K��p#�ǿ�Yu�Xz{�V�q�鈝����� N,� ���Z������qlh�qlh)qLLz�B���M�U�zh��r���^~�.:ox,|	Q�o/:VW��9YTӁ��5�d���7�{o5��4�q6$��O�S��Q��y�+�s"!:�M<'��IV�v�
�89�W�j���M"��l�g�]W�7~,���k��caCi�XK��e��G��(-ۚ��7D�[g�����BH�V���mы�۱|O�T�lk�����C��CoT��a|MC�L1��c�I�/�m��S�2�Vɻ�I!'�=Q9u��\M�\O�荢��,{Je���Z��9��h�Ɨ!e�mߝ��"zx���r�΢�4x|:�XŸìzG��۸t��C�}��eI{�gv�T��Ғ:G��$����V�b)��f'�҇��+�x�#v�+	����?Mv��cS�2����a�v�nP���)�Ùa���&μ��"kz��W=kEiR1�եj�W���r�Ƀt7m�Z$Hb4�*��L��d��h��'��މT�hqb��.��w$D��6�!�,W��l^: ���5��(B�¿�/��/U��~�[V�����q�Sُ�H��bx��	�%�ı�KC��?��͍���q��ޛ9j�M��� � 
o�/l�ޕb���1�o�,�)���[v֧�������y���{�����!��}�#���$u�j��� n�JG�XҲ�xa���]��Ŏ�|:�f����
�-k�F�H�e͢��lVjͰG��eZ�7�!�F���u]),*4wPXq�$1�w�d���d��C&Rx�ټ<H��������JD������~V��� {Ѷي�&i@;)'L4��'\��S��X4z;��E�o_�irz���]��Ƙ��2k)����=�F�E��NG�'�Bu��5��� K��i7�hAx��e<��]�Ѝ�]P�Z@�kp�8?��	f��[iEUi�-J���r�e���b{��-}�5U֮�*H��-/;$]7��ftBQoU��Ŧ��/�A[?��A<��w
:��5[���,�y[����߾���Lt}�Qg�&<{��^,Ì��H̥���:�G���h���g2�l��HUz�Ʀ�����tM��l��1�������m��ClB����g��_�<�h�ld��_(t�y����?�����?O��v�D��b?ZQ�G������Y]dB�u�m��
n�W;�t,(�!,ٕ�I{hh�,oV-7DW�}+�O�,�$kk�cD0���ϋ�k�C��.t5��b<�}*s0�+2.��Ȟwo@m�"u�����f���&�%u#�;{��C b����w
�J}����:�-�TW��)��zP7�!���i`0�:j,=x���r����<��f�J�\YIQ7˶Prp�7d4��q��18�/1���	���5�"}��Rˁ|�^���}�UI����{m_�̆1�q炌�!�����Ҹ�U��&����]^��HT�[HR����^*�B&a��}Sϙ wJH�^fwɩ?�k8�]zU��_p�Ύ�q�:�ªz���Δ�%�6��A���j3Tl�fk=(Ů��{��+�m0#��'@��@��~4>��b`W!p��44*U��]��ʭu��L��8���^���$b�U�{�wuL����bk�W�a�J'��փ>f��ox��d"���-�xk;��Q~���)"��;��ZO��O[����a����j���D��yYz�j�����a�����U\H%ٯ�B,7��:#擭\���,z�b�;]���X��2�\֐�^n�Zs�ϽM\W ��Aʺ�u��J���*�/m�,�&1�}=	�CB�$���t������zɩ���*ztCk��b�2�M���R�`���nr2�͏a�`V_�:'ȏ=��c���)+�ލ�>�����d�����oZ)���⴦����w���F'�1b�/��Px��}yf�˗��v�Y{��(�񄴞�����7Y�Fo��q��J�7��*@9�;槓x�(�2V��f��Blg����7�t4��S�L�`��W���z	��^�ItT���=+�Y�֪*R#J�xiq�ۦ�/� i�G&�u2{��Lk��X�^��8�^f��Y�JR������m}~+��)h� �����88��bL���o��|���k-	J ��hL�T�t]��-G,���&x�.�|(�tLYܵY���5Tm�}��[��M��PA�ѱs��[�P{*��ڀ�	�t߿��?��qet�x������U�'��5vwKZ�`�r�ߚ5hO]�8^/��ޗ��C�a���2N���T��(iUK��.����s�k#�s���(d���#����~��$��4��+sj�Q��.��z:�pn��Ҧ�ؾ5'ذ[bg�',A#��-�}�S�Ϧv���~	�PJ�Ω���=\u�p����J>ܴ��,wHwMz���|���Λ.vOd؛u����jiĻ�o^d�bU�Y�{q�R��`�5Zr�G���9o�R���d��ٕqC~����:}��<ɿ�L/�T?�p���'����<�U�VX<�Ix�U���Ӌ���������f�k��V��@��'����bG� v�����5�uzO�aU�_҃C�h�m�Q�E6���>)���}��$]q��C��5V��i�#�CD��4T+ʐ���WX�o�蛆�˻��-�^�m�T� ۲Us���`�1�4^Q�ω)��
.(.ê��7X�����j���iT�TD�2^!����w]nP��w����F"�;�mb�+UxAt��^>]�S������p�� "�|��徆f_�p砥|����W����ݲ���������o�ntDZ��1��P�c	��񜙑��W�q6=u�//-��Z��3��+�X��zх~Y�l)��mt�ӭ,p����go�m�\úx�~,d��8���ܧd���|����J�������by����u�(��NS�e:p��L�6^S�����8nӷ��Gq>ko�������l.��!Ճ�`&}��Z;�G]�v�6�����N�l'g�_'Y����@V�B>��d�������)+u|�$��U�Π��$}	�;�8��Ek��xiX6PŊ��G*ҝ�V��x����\a���}�n���G����!]��P�;]�ݗ0�;�wN�t���M�gW��p5�V.Jg�m>8�8�U�j�`�r�	���%W�O�K�?����8`��R�>�ΦП�uկ�\��;1�r���9��s:j�������_���>��؟�-�����~��Ƿ�?��?.����IГ򤗬)���) V��}Rz�+��v:ⷦ�_xE�yx�?�zu�
hi
��E��o���z�C ���WQW#T��q�S��"u`)��2!�9��&�������|Q�(�P%�|��@����z^�I���RR!�^���z?Ji<�-�^+�6g=��I2B���C�Go�R����3>�����5P�vW���;V��\3I߅V�9sk]���9=�dG3f(%�ہ$k�7)��3�J��(��'�M�I�O�y�Ů�[�Έ3�=EڻZ�X2��n�R���B�L�}����(��Ĳbs8��b�<E���Z�Y$��ZB#��Oߑ���?>-i��"�S?�X�|G��ɬ�#��2���8nK�<���x���%�}G \��<"�/�7M�/��p�?Y�'�����@��K�:K+W˽uHQ�b~���½���Ӯ���<Ղ��%4��4<t_��z�������C���5�8��}l~�e��G�;/ڸ���͠���ӂ�䊾E�(�>���;Un�}rW12�h��'��ј>Y`Ӗ�~��n�ñ�>�(��r;��O����7i�]7*6�U���+�X+1W���Ǘd`Q�y�{���.W�0Ao�#ݑ֒���fc6_[F�kɷ��K�A�с�Ȫ�U�;e��̊�1���ΑB��710'#���[�Z���tL���L�1���ߌc�T��c�Q��O��_KR�y~}��
�/����]�=�=$B���`�6�;�����w������ۉ�~��~�����}��&�
EǙ2��p�\Ϻ�6E�"ن�,����'�����e�� �u]5疭ǖ���*�Җ�ˇ�m�`�҉e��C Q�;���$}��親Z(�/E1r�a�w�{skˮu�t����]T�LY�k$���5Iؽ�7�n���e�:cKY����[�ò��t/��eT�|=���}ʯs��e$���O��3M??W;F�?_��W������V��dx����
��?����:5T,����-����
��
��j�&�s^�����x��e�� M�y�{y���k����E�yz����������B;�#�����ͳ��i"�����O}P2������l��؅�����?�a-�s;�z*�-He�"悛m:���?�8��=�<�방��S|Cp�A��-}zc`�_��S�d�cK [�L/?�=ݍM3����n-�6�1a��Xs��_�E�ֽ�(|��5��Uz*I-�_�16:Yۥ�:i��ߋ\<Y���Pd��G���$�O&�눆�a�2�PO��k:�K�}������� ����T�)�� ����������c�WNjg��j��D�\�m�?��ʃ^�3�ݮ^\�>-1�}�PX.�.6�w�=1iP��e��}+���_ђ ��\�e�YHw�BaN���U�����S�d=�؟~$�-NN4Y� ����nӚo��g��pgc���A|���|����9���?`׳[i�a:���~�*�ҋT/%�/G�=F$*H��-=���dR[��e?�zH��E�.���;�/IG�ނXV`)8�I�8�C�T�k�pQ��t�����k�FFo��H��H�*�ٗP*��@�~{��s;7�H� ���x�	�?�2xlǧ"��w/�.t������P{>���STvA��{���'������p�0^I�8����&s����'�!q���FnM���6�%Ѭ�U����t�V��&�O�!�:ؕh}�߳��"� ��M��:�<+��y(	7��v�ŰqG��=(��7�U�[�5B-�=F��/�\ȫ� 8��Hj[��� zI��gb�]����8�i~�L�b%P���F�ܞ�L�����B�9�q��5!ֲQ1�W�UY��^����]E�n:�i=	�<RO���A�|2�%VM]	�hGk
��c��n�K6P�	���f3�FO�tj�q�Ԧ9n���EN�����j���M!S�F��6�)�\Y�?o��`�4��2:������m-JtK�ݴ\�a,Z~�22��[U�E�]��ٱ��sh]|���]����\gu�)����m���ౡ
;�/ho���W]qy� �t�V����eP��S&�"G�z���zG��*Զ�uG�	��	�o������ݰ;���=k�1����n�
�r������Ud�}�x"��+�(˘����)Xg�1�I�������^>����Ѹ��Ч#��t,Ã�30�,�[4���(�g� ���  6���̗��f0������f�[o~{K�;. ��j�֋�7f�92q�C�����?�'�W+�����2V$�����@�u1~x�@ �ײ��F�������Y�"��<�E�YS&�WG[ݘ����?�V�x)�@�W�=�M���z���5jS<Hհ{nپ��<F��r�b�|p��eR��D,jߠ}���(;��]3��[o՘q�m�S��ڒI"�m��k���
1r3�hS�>�i]��:�ʠ�ȐB�+�f�q��t}8���%)uT��8�����T=��Ȉ�W�u�#�ӳ��;-cxM�1�kz��H��j	.�
	���ܟ��.�7K-h�R
���.,e/9o5uV��͸�
5#ݚ�����Խћl��5���b� �X����|��C�j%t%�֪�7�S��+A<�f�v<J�@�f�@S�^z᫼��p����ǎ��Z��Z�/�Ċ��7	���I�Q��Nx\����Y�,B8[κ�~�v��m*�h�.2�sMx��]�={]3	�`.��a)�d��x��A�DI�+.|)�n���&�[�^/s�U�;u�6*�Q�L�Ƨ��/G)x8�S�v�_U��(�5�46��roS:
$W�����Mnr\W�d�?~��SK�)�W^��w�J0�"�E�-���js��y������b���k:W���IUR�1��8��z���/��:a��P��P��)��e�畢��9�no���k1�r��$}k��Me�������Я"A�֨B����p���E�=�[dSI�2�������j��ԟ�X
yarJ.���h+��!1�$�j�1ε;P*.Ђ̩WIaD2DM��_G�d|v-�޼b�D�2��h��d?ҴB�֤!�v�D3M��U,�㈀�	��oy�~�a�����Cg��~6�T�a;�D�6Hz�0���x�תM�ܸ��I��5-�N*�K�\*�*��2���ݸ�V�NL�$@da�j�2A��O�[5�of���j�ZZvWD�u�
.��%@'6�vps��Bm���	�}���ar�6J�6�"ݞ�R�"M�Ӊ�
�	%���,�Ơ�[���Xdao�-�B��Fd���� }F�þ[@�[9K�6���g�-�^�Қ�� �B�,M�_\����[xZ~\�+���3X��F�F>'A�H��E�e��\���m3BӄW��F.w�)\�ւ͊���pV�0~jz??'
V o���:��P��5W_T&�*�u*@�S��mQ\.\<�-q%뇁VѢ��pj��|!��!Z��]��{θ��U����g$X|N�$�s�ۤ�s�6��R��>(.�#4�%*U??�Hn���d+�aC��v���q�v+�tkFOY$���嬉�L&�%�g{�n�0�`��L��B�'>ǞO�»{�.��5�[cZf%�_P��r9*>犤U��^1i��v�ό��ڛSb��
��q����3�t\0��{�BJ�5���(ֹ׺<g�� 8\�6�/6{1j<к>��o�]oۣ��j�5��Ϗt7I�d�(<k�ws������k�v"m_�D*�����#���Kf���PㄲJN����v�Q��m��@�[?0�5�뭕v�E�`�$����Bk��&L�3��⥼Ū6sOwc�q��8�s����0��&t̺tq��e���o��b�FhkK�� �Q��q�"�
��,�5���|���j��4ďp�xzfH���[
�o%P�w������8�­S��V������-��:p��E`�}���Xr
�'�ix�&���h�>-�m	�;���=89��h��DT�&d=SUy:ţΎ�}�î�7N��)�-oǅ��
���Z�N�h�U3�Al?�Bo3��7�~(6�aı�t".��n�+gA�`��\O$2º�vlz]���j_J���.��N�+�D{H�4�
SSݫ5_��V�W�^N�D�G"�7e@��R�KG�_�y�}Y���O���sԇ�}��￹0�� ������2��� ��W��'_� � ����� ���?=�Gi�'����ƜbG��ekQ����6�X���T�w�M���B���߷'�L��n�0�R�c�}褸FR��՝L�����K/ڨ�u���q)S��(g�{�P�� �y��ƵV����T��׭QI!%+D!���(�V槬�M6����	qq����{s�}�?�K}>������G�}��|��y���}^�L�հ#�Ҭ�[�;i��������b�B�g\���E�v:����K�Mń�-�+�u��=��;c%ܴc���.����9'�gp3@k��b��S���ҪS�
V9�*�o*��2���_w�߇����D�$}9�\4�D�U���>_�u�����򪀱��V|��"�_�6MNv8ݞ�+s0(~��;��3�%U�WQ�Y�R���~�b�t��=%ʑ#�H_u�wF+s�yɺg���.�Ƣ^�]�fq����1��S��?Ιۺ�k��>���Da�UB�DO���U��v��۱$�<�-ہ��Udx�"r7y���W��[�p��7��мs!�1G5�jf�3�:��Ki��7=�`LYȫ�B����OaZ"j�U�i���̳N�~'e+�q��y���k��u۲U���c��Y�m7t|��wl�js]Dt���71�!�
݉���c}�s����#[*?dxSs��:<���k0�_六е-v{�O�
[��8&���S�[?*y�ʣ{�KY��r���C&��H��[I�7�G�M�]~YW���N��]k1`fR�>-Ѫ��KRVM��޺߬�t��>̡���i�&f��R�0A�:�e6-Ѷ��R�nh��ax�Y��Q ��QI��O� SZ|�O��&ІX��$J��S=#ӟ��/w�Iѩ@�ˁ��>�~����vU���Jڔ_g��e��9���k&���	�[���7S^�B��V̾�x�[9�?�˪A;_X�Ҙ	o�:5�g�g�������o�=�i6��*b9]$�{?�ʛi5��Mj\=�-#[�<6�FaV�s��ɠ�-1��JT_t��Ҹwh�e�A���l��d�9j�%E���E79<ym�N[&6��-��yOy���u_�P�����r�	u��&���v퍎�;Q?���68���������jS��v��<{#�2R
/�^�`����*���}���-I����U�������-����R��8�-z'���|��N��ڝ$��i_�n�pl�/*F\߮�T����$�yf��<E�6T��6:^E�r��
�d��~@F�,�U^Oι=φJ����R�}X=��b]��a �����'�^<v��}&�ݥp�Τ�\;B�����Z�>������ݪ�J⮽���p��Ec]G��(]����:5��=����Mg�3ع�������֜}u���7��CR��ҫ[Dn����ܼ����&�p�Ӽ�y�\��@f�����^5��>��&��^�5���Z��h��^��;.R��F̋���},��c].F}v������(�,b����:�.qdg��y8N���j�sC����S�ß��+?�H*����O��G���Y-]P@���Z_����=�Ťj1k�A?�1M5vW�@�\v�>[�����6F��!�S�JYs{?�	���g�*nq�3G*�xo|<�fƐ��T#M�Wx���N��'�)��a)?��h��j�i���,��Q����!吶��a)_�1к������_�����a��w1�����J ���Q�e>:+D9'k�w!�pH" v"�3�f�P���&�-��R4hs^�)��A��SH��p��d�C�P�.�j�jqE�U�6����� ����!އE�q]>�<�z�n��.����X���ڞ��_��7�a�)���iE�qI�7�F|}���dHU��	���C`�	�u�����J�0*T-z$_[���U��WV�Mj]R'ކ����x�N���hn �Q�E��Ob+�/����.=V_�˵�x�2d���[�W�,�X9!�����R��t�"�zH�QvkϷ�	���/X��7b[���Z_�a��MyV/@|s�u�/�����Ϭ�ah�W{���*�5�dˢ5�r4B�ne�I_զ��H�':}�葂��Buќ�v���U��tF�J��n�gV_sM�0��m�g9� ?�n5֍Mc�g�'pI�LDi�`�m��f����}��U���0���G;���s�a|����{��n&�F֢V�^���:��t����ڵœ��y'&�'����bE��ۿn�U�����2�<*�������`f:�V��c�?&\�5��o��:V�N���]#����j@8��ѻ���1?�|m��v]8E�WM���~z߇����A?��Ժ�h�cP�*���L���\�v��{����hº�
"�v��/��T��:�|�z�v;�vZj�����l�z��Ԋn�+UW�ߩ?%���}=���tD;Pܗ_l�v\�˪���,��F,u8g�h��9��x�vBL�/[C	��k�態�6�2P���4�D�t#�d�0x��2��ه
5��7�_��ۺ<㘋��d��%&3U��\�ƒ~cn�Q6Z%ۍ�����_d��T���U9��r ����O����j����岨nx���ڜ�"�}�ݴ����YR[ޱ&�	T�͎�����P�$�??`�̲��r���ܪ{�b�5��F5L��ZP+�"�MǺ��4������Yh܃q�p��Y�ՐUW��k�߱�lj���wktg�_�x2-Z���0�hz ��Ǣ׮$�|[܃��MN���(ay�Ln<��J�o]��Kc���nd[c��aV�άe�x3�4#���o�kΗ��g<�I3jw����{�[կ5����b��}Z[��ҁ�r�K���z��*-��|໅�J5��EO�j�M.7Jr�lGa�"�E�
p^*t���F4���u>�b�Bih|�K�����/�l�֋]:�s���J�%�:^���n��ى<I�.����sȥz��2�y`c�?_c06!KwkMع �!=�贒��G�(ԗ~z]ic;jc�.����A�5���_^���=s�I-��>��M�Nt���5G���P�\)��Y�I��ى�կM
�4k\t�%�����E��S��.�O��E߫>ߥ��58�N۠�c�!���K��4[A�A<"O�{*�PD�F�/RAy<��W�w#�l;!l���㯪��l�T	�ƚcb�~�Ҭ߲�Q/�)	
l�ZxД,_�f#&Nd�z޺������]k���Kr\�8���(ў-ẀZ���VL�G�苊�aL����q��_$+Vw��х}ۣ\��ӈ���-����dV����n�A�][z�쫧�9W�C��`]Ӥ��ZRڴD�$��u�����yM5��R�s��<�`��O�Q��
��y���"��	���i �</9���H#��eR�RjG$GjW���\�١��7{�!��;l�F�*(		�[���K8��w6��*��뎽g1Z�\��c���k�U�Q���y�w��P�e���Se�Fٳ֫��ҩx��x��ܺ�h����|b{�U,�D�̙W8���s��Ҟ6�O�/��Y����[�f��֎�93Ȗ�)�w�����O�q��OI�����L�Z�f`U��z�~a�v����lʵM�_��a��l�en|<P��ӆk~����ri@��ۼ?�btH��,9ڞܕ��m1��ˮ����%\~��H��=�M����8-{���@~aE���s-3헶~6I/
Z�aRV����S�������XWPH1�;)SRu�������}ع/�\��'L��科5��K����j�|�>|kg��%����=Ί������Eg�>Z�k��X��Ҏ�����m,]�d�M�c�1"p%�lӽz�6���_C\k�c�����l�]ת�CZ��h6b��7�a!a:����oK�T�4}�s+�Y�kr$$YwI�[3�7�/��|�&g2���Jp�0W�����>PX���^�Lk��>Wk���!����jݝL�|�z���&��uwBow��g���9*ȋq?��0�%��3+��%��&R��f�[rW%[���a_t��\�F�P���5^�W��\�����.��*A_0']Wy�Gw4���GI���Q�V��-Y"�
�ԏ��X�&.��j_X�w���v�^G_�*L��x�0:կh�*���o����2u�^�����C!���O�;�y�Y�b�&�� O�ݬ���Ha�+Ьm��d���Ʒ�7���v���aMr���5�X��Iއ����\�xb�w+��*���̭�cgA���3�M|���}��Ĩ;D�|����vn0=y����p|���*��Л\������s��|�Wj�0c��_�ZqU��=Ca�μ�p���k�]��ΪJ�6��I�Ͱ(��_�O4��'4�n:�9u�mK�w�7wF옅�����5�dg��g�F4�3�T�5�d��,�2�����O1;Nm�#\q��aCu8��M�-�>n���@tK�}>GuT_���e	������H?�����bݧ��hK���(aZ��&��[���q����DZ_�^��L�O�iD�֢���:�������w_v�Ɲ˟h���S����j��v����]�}�eM���1��h�57��啝����oϰ_:s������a�����N���s2���K<���fY�k�nA�@1m- j�E����64*5�u��U�D�s�}��1<W�0,��Ws)y~�)?�a�n�bՆڎ����02��׳��z�:�y������4^��_��f���^��ϴ�%�r�2*YTIZY�E�oV��۱u�r��|YtG��������jyEϊ����4�3��6�;�Q9�,��3 �V��)e\%":�� '��f�޴IT��s���9�c��n�a��ϯh��|���?~���nKUZ�Ǡ�ڇ�u�OY?w�^q����~dL����MU�hG/���d+���y(�����c�o��򷶪�"���=.Tg혝������͆�re��O����D�/4y+��]���io7V�U�v�a�ڿ�m�^��R�]wR\�EZ�?�rC�Z.P�<:�)秤SҲw�?c���!>st!�}v�gkG�u��'��h�e�S�tg��*E��VYk�᫣Wؼ��xOF쥌�M�1ƹ��2A�H{�iś[;��S��qO�"U�'���*�m�Rl,�wſ
����̾V�vV,IE�`>�c�Ò�8�v��-�<���1
��Bd�]��;�~�5u��V��̊cO��:s�"�����O���/M�9��;*����QJqt.6a������/�Ѝ!�g�����1?]���ܑ�-�3���<J�㕅N�c�|{�$�W���]�u��0w�/������Xcy��Ă?�.���3`�>N���q�%��\�[lŬ89�4���Q<��,�rr}��f��p㍘�l\��܌������p�*ά�lo�<w��k7�-^���;��s�4��қ�l��/舻Ŏ���lK��\��p�eAl�֦���m�~�͏\�aQ�[܍��k�K����p:�n؏��g��J����ٍJ�h0ϙFq��>���-,� ]��EX��Lq��������ye�obj[��[�V,���ŎNG9n	��-Lݾ�J_�o���5E�/�=U�������[�/��j��n��i8F�6W�[M6�jZu�;O�+�&"��Yd`d������}vPچ��?�:;�b*�m��}59��㶮�n�.�J������<]�����K�B�9&i��
��E�aƉ����B|�oxu�>ONF\wqPi�η=�W{�x�[d�������d�^�D���Yvzf:�X��'衁|7Q�^�W�Ғ7y7-go�yp�����-Qt"���q��.�;������-2�V��s��.
	�t��K�D->ؿ�U1E��^ڝ(�.	>)�g�dK���8ʜ��/ݟ�w�����H��	�*���i"p[�;�IAJ+���CV��{������~�����-�4{��5UQ��&���X:~�9]]�̹잲v��s��3
�ʺʙ�iW�6���u��u�w�s0��m��)�R6ӗ�L��?�����ƪk�}@��6�Ώ�J�dbPv�nޜ��/(s�r�Z�|D�r��Er�g���s�f��sY�Y�8�b���HC�(|���(�5�?;�u�Y�熯��)Vul�ᴊ��k�Y����XSgn!ׇ?x��4��N���kF0�2%=T�r�η��:Y���d�E+%��`�IS����y�ޒ�9��E��42s�z�������R�m��r�(�Mb�I>lN���Ke|� Ϻ�$D�b#R�!���D0��+�`�x@z���OXN^d?��������^��?�_�֘ꫡz�����_�I.&�S}�η�@�y��vv�����aS?���6�n"�k��t�wO�׮w�P�y]5c&�P�T�z�7��
/m9f��[f�~�/�;Z��ۺԺ6�ԭ!��킊+q\�r����[�߲|T�׿��;��N��LK�ʹߺ��3��J�tS:���������m ���
'ij�y�}#O2�*kVC���k�Cj��-fA�q1?g���Q���Y��'6\�ҷ]���̰_
q7�+��:����(��Q%[�13�H�M���3��٦����ЋJ�Ʊ�.&>q��������ܦ�����,v��\�i��`�����xU�c_���O,?����6�5l�W7u-@7�;�x�����҂�7�l32������|�g�f�Ǚ��9'pa�k�o᪛
�x��3.�`+��f�ጘG�G�~M��G/r�>ېJz{���خ�6'�/F�����b�+�Xh\�������&���$��_�y?���g�����Z!�bv��e�o3y�ػ�?j{��N���}��*/]�Z��)��qᥒI��i�0�pu��>l��D��X�t]r��ܛ��,\uW,����)�\j�Z�}�Ao�[�ב��7\j�mk4��dX��[���8j��U�]�5t�6��@�a�W;�|�c:k$>�
9\���`K���>�y�a��c��7�e�+�d&d<�=htgf��W�T�l��k���؊gx�1"�rؘv�e?����:	�m�@���(_���Cv�����粦c޽Lĵ\���x+�l���L�cN�Rz,�¸�c�Ո#�\Q���X���.���k�%c26���Y�YI��<�/N9v����\@��эcci�5[-�c�W��ȅ�m?���\6�v��s+���$\��6t�>�67)R-�ʉv3�|���ry��m�_Үk�(����^`x��ڜ s^��p�������S���Yj���z�<i�3��Cټy�$֨��.lGL�\w)��Rإ��L�n,��~�<ʔ��p��;�b��&��:a϶�6#�`:���9VW*uI�����o�t���W9���j���
o/�*3�Z��7_��f��I�TQw}q����fl?��;�5M�~^�2��z ta8�t/8'��n�(vS`�&4�ت�|�*7�mnh��h�d���X���9t��ֈ��7åϲ��@_���j��Ω�����B�j�.uN��cn;Ud�JE�5��vt�Wy�Mg$�g*<�ߐ2�nq3�`j��Y�*co-WdD���,Ǌ�E���#��#�w��`� �k���W�ys_��>�Q�⋻d��p�ݳ9]��5�����*��"�@�ت;(Ve;n�t���t`	)nӹ�7�j��9;��@N��Y���֧6�U��h_g��F􄹭��9�ĥg�tWc$���ո^r,�`��Rsz`^u�&��\�&Ϗ�ޖo�Fdn%��0�f͠��?�)��启���_Z��\�~~����ּ��ˍj�M�R8�~Z9��Rc��\�t���jn]�Li��k�ʍ�Ɖغ��o;��T\�s,�p]T��6�Lr�=�6�=���?�T�D�v�{�4�\[+W��.��buݰ�������|_v�����d���y���s��'���_��T4�O��-[��q�6+�z6ĥ5�XW5Mg v7����z�}��:)�䔬Ր�����sq_#�j��B�+��i�.J&����USv�"8���G󜒮����_����`֭u���ۑ���C|�FgRD�C���8��}y)z���GoN��YZ#��TB��s�Pej����}پ�Qn9�L����a�k��8̌J�s����آ%}��>��FHC���5�s���"ΞR�L_ݸ	������m�v-)�/��?�|�ʖ{&��{��:�=b��ᰩ���p#�Y���Ѷ�Y[�s����ەLMM��펩�/�a#��w5�rn�71#L�V
�D��X3�ix��BT�.�N\Q�L�%q���	���ɢ��:��֖���:�I���!!�JI�����?y3�u^;�@$�{ʤ����J��+X�du�ل��Q�N���k�;�����7bL��[�ۄ���]��O��B�k�7�r�5O�o����z�KU�V\��g����� �4sc,�I��^�M�sK��Y+͵!��\�F)�nE�3m��2���p��q+w����&t�yAXvzI�PNj�V��hA#oT�VyyX�5W;��V�ҋ�.��g��v�h�\�ug��t����w�7h�|�։'�����ʭ�6����KO4���͋Ag႗F������-���F��Ԟ�fi_��U�߮��ן�-�/y��>fOV�v��T��5�2��$B��Yd7g-��z+�|��CLH�\�ꜝ��.[�{�y9�V6� ����.k9��Ou;{h��K�R��	i�q����J>���|N�m�_��p�p�����5����#~�7���Z����@��:~G�Zõ �����}��Zo�ֻ�����9�d[���;Mk]g�K�'$ziBS���r>�aU�P�h�;w�\ئg)F��N�ɐ�/�U$���	�q���"K�A��HI
ՍL$<�ׇU����
��Cz�-��������y"�%YB��N<a�9��d�My��{Y9�f)���IW��w���#�&B6=�,�*)�����gV�V������]�ض
���"M
���+�qhl A�q�G�o^鞖pi���߇��֬��u�N1�5[*��5�#���+3(�Q6����յ��׹Y�mXsJS��z/J��J�lZu��K������K:��Xɋ;�}���͝��G��t'so�7��u�R��i�EC�͈_O�;�h�4D��mk�q<�v:9��a$qq��7��B�.U��4̠�"�jw5h�a�DmĪX���{��\�T�aM�U{g�DY������;NH��^���VϷ�c��+X����)ϻo:Wk�R��`ˋ�c9:�Iި��Xf��.�n.����6��W��M��)4�-�*��2GT�P^J\���~���b��/��쀕����<�]��YZ)��i����t��@U7��ޞ�$љ���:W��}w;i�йm�% ���|�_{v���n/}+z`u3���.օA[�nf�\{��@���(�2���z5wz/CT��B��P��֛�д.�w{��߷.��Z�b^!�݇���Ax�u�_���ڇC��	���68�ܞ����ko��fB&xv �X��-�.uf�@��w�ݲ/?���r�e
�;�}���;�w���s��S��0��?�g�o8�q�p�)NĮ1'fp⤕���f��$AMk�[�t�`7�،�M�:�;A��#�'G�a�bV�s�����<��*FvuhT���嶖t¾�j=��]:�~�0�J%B�K��q�P)�ߚ�Po�K\,���u_�އA���˿\-�
�����7����D��1t����Y��W"��F@"�=�Y#!T�;�û?�D��S�Ij������j��h�T1Z1����3�n��Ų��{�f���n9��e���(�9�-��QNJ�7v���˾e_��ƌep���=l����u8p<���s�C}V�޶���z�\z{a�KZ�ci��#��8�mf��O�!��!�F�r�܌��r�;vmT8���%��-6(�@g��\�@���RO�^���]`�rw�6ʗZ�����ҹ4���e�Z�3�].L��/��`�WD��b�n�~�c�IۇuXC�:|{[�4�#3�Y&a�n��m;u�U\~��G��f�S�6
v����4����_���K���s��K(Kdǥ�{1*[2��):��ʌ\�SE�:���0B"�����e1п4����͐�M<��N��8�X�rI��7�I�iA�s�ˎ�z|1��0�=F>Fu�]\�\���� 3����݌�%�7	��b,�݀��m�jC]�+�J��;:�7�@�'b>ۑ�9�Pף�U���;�2��y�+��0ݎ|w��;(ӪyX�G��i!�����̸��8��qlt�	����0�I��(��+���N������>��e��B#4`��~����Hg�+��%f�C���-�\k��Q\.�s��F;8�ʉN�h��3���A���=q{̃NL�C����_�ڲ)�K�~�����c�Vd@���~�B�t�^T�N��ɐ�����%9�L�K�s�YB�{�`H��������dx���yḅ�� �a�P��x�y��`�N]5s���Ѵ��ӡ]�������]��~I�h��pj{zw�3l]���K��썕M۵Ř��|[��\o��a�b�V2��61_�^+�����rd�1f}�Ҷ(��}XyĀz��F�<p��fE�m�o�b�ٚ���;�T�aJcNd�������<j�7����,;D��I�,5{��or��Z����c��J2n�a)sn5-v�My�6����=�N�g��A�ЇN-̈́���}<��W	�y�h�*HE�>�+M���[��OD�"�?�	�e�!��Ϯx�&c�3l��{�鴕��2����U'
-�o�	T�+c�N[Fޖ�gb���=:����0�D��ntC;�/A
y	q����O��s�p'�Knp�܀n+G@�:(\9�]R	*T�$�w^�\D6`�}G��-�-]?�|!�"�;I|�~�S������D�$����<�'ӱ�}G7�� �m��=
~�l8^���=�o��D�[H�=yzr�P2���U�eh�����B	H$���pv΃�o�:�%�|���g=��(���g_{I��QV��y�y&A��Q��)����t���ϙ��p�&eOq6�t-��%��!�@��,Љ�
�>P��Dr��qM��c���Q�>��9_D"��
�7���2�����h�o��w!s+b�ԧ�|60�G'S�mRh���U�P�'u�B3�Z��T���xɖȋRq#7�1^�M%��0�D��Kt����)��8$��m���"7�ѳ�{z�B3L_@�)ZxU9��P���=��g��;�4l�.���'��U�2 ,	DX�o����{o���K ��~مzP-�����w��w�ɗC	���ꏀ;�M!����!zb��)�)�:�V��K-����?�_��$���'z.�q#���彿@���5��F�S�.���u����=�u�a�)uhx2aO��dG�A[C�+�L�W1�:#A�ے;�!l�}z�{ ����P3~y���?')r!� ��#��gA�S�^�aH���Ƞ�:��F�L��p�	{3�p�X�D��B�#�>���|���xl`�����dN//ï�Z�x���v��h�T��mIG
�>t���ꏬ�zl@�y��X7i���;���0�tr@����M�9_b(����M�x�ϻ0}Px�(��^�)()��9�l]����9�iK:�AV�w߁�wޟ���7a���|I]���4����xހ�~����ߤ�� _O7b�JǪX�܎b����)�&����#v����d�Up���P.��# �k}O��k}}�?�&����p��������K3�S !zb�!.�3d�xQ�>����]2�
�=T �P(�!v.K仁��%/��@�\�,�m=��ui���zI,s�;������o�s�/�!�59՟)`uG[8�d|���9?O���ȟl8}aI���ZO��^�
�*T��/�/@�t؀�#I}2,E�v��9�R�^���h@z��I?���xE����╂c����G�>��黰NTTZ���:�=n�jXvٗu�kK���Nh"�Ɂ���o�r����Z��2� �d��`��x&7Eb����f_~%J� �&���'�����CeS
�&�(���@��Y��S�qD�^},l=j��U$ZߕA
��uL\��̋�� �@��B��Dh��RI 1�\Y9��@n7�4P��&�À��\��.^�*��{ � �!��?�)��B��(p'���a ��U� �������*)��	�u���S ]�ʾ��X�Xe]M�ގ���d}詖���h^��C����H���&���J�Đ�B()�C�c��20u����0�>�:����o��\�#"�]�S�z{{�Xt� E�_F2?U��=Ӯ;��\W_'J�~u���s�u"Q:�/W	�����[��ʦPg"���`%���B����(<v~�c _�%/C�|x��r�uQ�,p��W�9D7��8,݂���>�>z���X���WX_BwG�-[��E����:�� 往:���X�i��4ó�4�K`6 �M���P]"�/�/�{�N`L��t 
i9R�����=��y�#����NF�@�')���|�����~%'���:�m�����A�����I�4�|�����Gɠ`Le�A&��K��JA�O�U%��D IY���=!Bz�:�܃u����hi����yn�A����E�0���{0�n���.̋X ���zcrG�1ۤt��{�a���i�w��0��??��K��
�~J�~؆����H����		��t��߽��-w'J�pa��p�~�)b��E&����O���ذ�ܰ&�M��qS	����-�G�%d�Mbn��m���4p��9I�����K��U���"�xy����'��$����B���4K�x��x�4��hJ�{�D/�߮/�ˬ��po	��f�Q$�.%�0P"Y^Ц��{X����Id��Ϻ'�H� K$��!�G	���Q� (�}�I	5sNS]��0�B�>���i_��*�[,�>>����V�qZ�pCt�ꙇѳ���7�z�$T$����$i#ٽӉ,����h�"eȺ��ꛒA�Ζ�`Qf?�3'�����9��'�

DD����ӊI���HD��G	���3y���h�;���X"�/��HJ�B�eG<8�Ch�4�&��P@�P��pl�|�%Xf� ��͖s�,�	c�D& Y$H3��Y%�(�P�g��Z�á]���`���<���o'2m$ ��G��"����LJD$S�� ��PNؑ�?X��&�C0��62Aq�4����E����i�B��X�(L2��a	��'�J�Wr����3P�_�T@{J#��~z��	:3��
~��H�k���H	��0%��;�2J�y:�4�;Hp"��"=���G��T((���� �x:��
��3����Л�	��"�RNI���o�0u(�ş���C����f
�)Dl�<�A�>���i'=����𐇆L�LzT ?H(5�1�����ˤ��Bȳ�8�Y���~P*"qJ�攧�A(�� aO&7����Z�o&�����G��I��@=$>���������x�P�������C�`)��񾢄R�{��H�R)��2�8P�m����1P*�gE�3큇`�" �l@7�(a$�m)06�)�C&D)&@�œ�3z�	s���"I�(=� !�pAr&	(J	w��;`qJ�<�p�?G@���A��a(0e0�0)Ј�D���#�y�,��lA��l�	I�D5��J�
t�_�a��dc�?�W$��?X{"�p-%X�RN! ��Q��%P�BJ	GAP�
Y
ҁ��ý����$�f�{"� ��FR<#HU�_�=>���ɫ|���Zs�p�0,���H�¡�K��%������ƆH�)g#O
t�<�@Ix:��Fx:X�� Qe��@�& .�W!�k�����JI9:�pq**U�1��r+�'qIa�A� q�f���� ���9���0";���*0#�0!ɐ�A,��=�@�����<5��Ѓ`S$`/2`����9�ŁL�*A� %P�E�ix�
t�&�� 7�?��a�|R8#=@CpOi"���Bl08�!w�9��?:Mb�x*��@�G y�"��� �cc9JeL�
�҇
:��0��$j�
���.���vӢ�/��k!�\�q�.Bz:�-Pw�0�!b&� -���D�j�J/�(@��=Ȍ�z �
�@7%� �0�
fD�"R2rM�T�I�{JI��S��硄��!~�2+tV���R�r�	#�8X�G���F���-�ā
0>�4�BI����N��c�	C����E��=�&��)�<L���Ya�	p�I��$���9�"A�(I}�P��k�(�1`n�'��~����)��MO��R�`���}�l��N������}>G�IB>G8�b5�oB�;cEԛ
܃�PW�� *@Ny�(�L����l�pPRaHy?E�W�Ui�a�D	X�)������G0�+
��K PB�s��ȳ�)э?H� f�'=Ԫ�H�L����7 +�BsK	T0�Y��3=�!��@|L������j�i����/����4����{`�(����a��C�x<�	H��@M �Ya�p@�ྠ FP�/^2D��y��qG��S�C��@�R&�gރT-�{�C<��J�z���??�y6�@͜>x�}��������w�
�[t)�'8��#H��I �i,]��6b�Y�Nýԁ� ����J��WA�1`܀xet�����"��oM �w}�q�$�{�n�P��R@Ft��\2%$u�i� ,oZ���yO�8_��eC�E N��"n���2U�%X�#>@+�W[��Ax���1����zR�x�$X	�V�<����� ���_3(d�4i��P�o�����vH g9��a��\bֿD�Lr ђ`D�'�W$���x�1@��(0@��<����7T0 ��,��"O�����X���A����A�+iT�R���������ZY�	�����o'�` �?x<.�ݢ<r��p�C&2gl��������EdK=H��bF�@�x�]	6VZ���D�o�f�O>V����mhyF	�c9GL���R���,��7�"x~��V�4�ea������BM�4�{j��C���?�bwNq=$�������<&�s"���%�0�A	���� $d�T�J�����QY�O�x"�f�uX�#�ҏ"�kD�������>p]u���PK   ��T`J�'�(  �)  /   images/1e039584-5af2-406d-af07-82deb6d77547.jpg�yeX���,www���NpwwKp'����%��wO� ᒽ���s�Z����鮪��y��u���"+)#	�@  z�� >1U	u%U^K3F'sKV&wWkKY)Ye	)���$���v�n�$$<,p�k� ������A�@AABB�AC��A�C@����GDBCADBE��G�BAE����D@�����A����;	��$,,"<"��7���0�#��� 0*�u  |��������@o|�q	�v����&�u@ �=�Fy;_M�� F���Ռ  ���ԙ}A:��� ���q ���6�S'T%b3]�
>�'�|I�w�%O�l_V�]F�<:�Դ�6T �e)B�A$p�ڜ�*�����H[�ދ�Ǝ���.���-�z+�|B���*&8�8����-G�������A��˫j_��=��T�F��y�y�j�S��k�~.�i2�,�ߺ�ؿ�;��UC���IDC(BD4�S���:V3̷4��}����'���?�y,�� ��;�:�Rѿd���a�I�(��<@���T���|�.ލ��#o�c)�U7����^��R��Ӕ˴t���9�"@���i(T�;�K��Zd�q�g��:;�/�<�Q��?|_��v��e;�Ԟ����O^�
 3`#Q�Ա�U�n�=b�;�8+~E#�W&zXR���ޒEJڝ?��;��-糏�#s�0�
��O5�����7�ľ���t�r\.��[����A	�����/��
~FC%�I�aI���<�իF:���VG;��V�Vk.v?>SĮq��'x�*N�8��nlF �7!�Ҳ�e<���k��f����CsC��"���/���Y�?��x8o֟&�(jT�7�����+��>1%�1�p�}����/�v�m���'��HR�\��E68�����G�l��^��r, Q��vE6���B<��FQ~�l4���'&����Л'0�  H	��*	��FE� �@�D���d�f�4"�z��!0o~��x�\W��M)3<�NU�?V�.m?�;���r7�;�T{���ݚ����|����=���e+.�y���m���0��ϛǗ4����Ⱥ��~��w j+���h�q	�6$��a�#��A�j��IH�S��p2���!X V[�S��̾�}�Y�!_G�fZI���=D[IŜ8|��D_V�%����d.�g����B4Iq;$	���c���՗���l?��>C�k@9f+D͘�^{��F�3JIؓU�P��fW��g��sk�+@Mʬ�V7g�!�~?�X"L��=���59��w�.�h����Hcک�tK�$2NC���"<ҽ���Eu���]%L��֠,�'�:#o�$<�9^�~2T��83}��N[#�>�l������I�m�9^�:8��.����L3=��4�{� ޑ�2Y�T�9c��k-�����A���={��@�IY��*��G�rB���~�JT<B��_\���m�p lD�fE��܇��ؽ�M������(�v�����eBSUw����	�'L�z�ѷ�Kw���Pf��P�Ind�R�%T�[a9.��7J�!K��=6�ȭnI�����Rٕ�^��;�CR��R�e���c	OhcP�3�K��a��+�AE8�1���4�چ|����#є}�d�kTZ2�sZ1v���Cj��ҭw��Ƙ��:��?3�C��F�J[�ny|�00I��ND���LΓ���X]����{����.������{A�	!w�����3[�7��}�S%-��+ú�Ə���E��Ӡ4���J5��G

g[��a����~$�@�veYv�*<Ӯ<�tiI<rlj&̮蹭T!�IzG�np�7��Dȵ�Bw�Kb��n�f.�f����K�Ky��s:���[ld�{FWғ;��af�g��Q�G�>�ε3Ջ�Uu#�5�Ѣ�=Iw��υr�֢H���S_�|��-��k�)�g��Ѫ�O{C`�_#[�{�*�����p��x��R��
����NW�`n����K�߽�q^�s�|n1 ��,�8^�f𰱾��ͻ[L�����Q��@�X��	��O�j�`�B���/,�f�C/�4}pz�S�
��B��ޕx��s����K�l~>V?�$&:��,��Evy�w��/c�K*�"ä��jk�7��B2�T��r�Ry��l����j�098�Φ&\_$�j5�O�Z6�
p�O}�o��'����PPYHHYE�!�	wo Bt��Ę�@�%P�ǰ_00Ȅ�ͅ�S]Pe�>�\ۅ?:<]x����&�ot%{��ox��o��6=+�:����?+@�]�A��N�&��)�x@�#%Fm��Gz��q��6��`y�Hj�	o��ouY�T(L�%i��T(\�����@�OU�P��tD�aTq����o���AA�@C����݀!Q�H��XE��P���b�'&}��!!gcW��¤�5q�X��f����?!���[�o��y�|\�g��-�ۊlur���)0.k��G�}��`�)]����S	{S����\gٌ��h�I3��@JS�+�9��
_�`��>M4��뮻�!Y��偼�۫ެi|�<�~i�3������N`r����{�8��ZKc�-�zR<�G���'?�-�h�N
�+>vz��gh���ܮ�Q^\�fyvta��� 6{,�o+_�pZ��9�J���EC:�i�2z��:ת �dc��L���w��m�B�>Ʈ��L���`�� �GC�,��捕���yI��2Rol�/�'׎�7ô�U��%����`���\_�Xz�;Qܷ~���~ն����=�O��*A�fuY-�����D&�%�.P)\%�W']��YR��b��y#�޹k!�^�%=�d����N�*b�t?��!�MЬ`�3���f׻��
��I�%T�~�����n�L�k���s���$1���8�ͪ�f�LϾ�����O�N��g��H-f��ÂC�����>�Tވ���c�8�I��L\i������{ƾ{�Y\�*-��Ŗ��O��=�v�|�/����Qa�Ujn��׭	�s�����W ����@���#`�u�\��@5�T�r�j%�r���q��:K�Θ�N1ـ�HG�xy�>zfd�5IS�Fҟ��ّrL&��{�P�-��y�B,�Y�Ad�,��S!I\S0}�5it����fd�^A~M�0l�ڱ�6�([��˻x�C󗛔~.ʣ��N�|<w���F9Ͷ�1QMwx9��;2h�h�,?ͷh͹��aQ��������*�rVW�칭%�A4��m��ʦ�\lLM=�����Y����J��lͽ��}z�F;����n
~�TR� e`�,��|�@�,X�ؽ������ېA��A�W�����~����Ÿl�GQ���]�MYy�i��}�]֍J�z�n�OP������JAG@�G��o����/���F�5�M��c�!�+�B�ne~a{��B��'����yLx�l}�*N�}����`l'�qSC�Z�r�:����p�H	�bB<���K
 ���V��l������Dm�	��5)��Kl���:(E|����oi��P'	F�����s&�B����ʶ��h������Jz�վ3	�����{�Wf!�������m��#�:_��%�}q�D�w��]�o�>Y
w�؉`p��5��Ό5=�@��j^3�M�"��ݷ�����h߁M������;�RI���Y�b�@��ʭ�ouI�t�s����b�1�K�@�
�lf�(���{���Z M�+,ggCz,|��K�HSb�yŕ3��0"[(��a~��j��r
��v6��`�h=T��d�Ll��򘺯d/��?��~�[���QZEV��sY^�X횫�:��s4��AYR�7k6s������MK�o������d��fN����<���u���4Jre���lLQ;_�0~�+Sm����P7���*��ťJ1*{tT3-��	#RK��ҷ�٘�L^�b���BmU�Pbߟ�
H�������*�GcuƗjܲ�Y!R<��N?CAk_QS�u��6� +��?(|�U��\FN��5�I�1�����)tI��e��?�Oa�&F�h���s��ȅ=ʙ� a>U�=g�U�V���� �1V�L����� )�+���,�@|٪°�uu�Q�$�e�ا��w
?�N�q6�4o>ɴ'
{l/���}�>8ػ�QQ�ޔ0�����G��nG7�Cg�w��z���	�䲝ס�-adML�12��VR���N/��7�Ȇm[�%�{2��~[��k5�����;��j�2��>�{���̃-R��0HTt��)�+���6^{�En�R�p��q:�ߥ�#OX����m���n��w.\��)�i�s�4ŇM\#���))�Z�Ŷ���W�qAUaGr+:mA�QDVt8���g-#b?�tF�� ���2wt�Y�(eF�H@���\��l�?3Ƽ!��.�|���>Ku��[-ׁ�%{4SԬ́���V>0�b�ւ�g��y�Zr{�����p�h��vZ��X3�,�.��B��_Z�+}�%�)�	�n_$J)�1�!����<$&�c�q���ճ��3�8ίhe���Т��݀���7�Ti@ �S1vN�Rw��;�m�r��dT����.j��(���$��ҧ�hu�uR�~*��"t�#��*Y��շ��2��6�3>T���("��.�Q:Ep�<�,bDg�O0m��c}N�M������� =�+H�������>]���)�&���~�����2R�-���;�H8D�.��j�z쀲闑`�Ğ*?y�O�r�h���|��l&�RI쉔�c���S���Xd*��|r���A����\��w�xDj�	S�:���G(�?����%�p��br�MV��}�}�-�Oy��޼��~Q�>��Z���Tm�W@j��!�Ȯ�2�J�ԌF9=�?��>C�[�Q���R���;�i�e����V�wJ=�q��8{D9郯S/&���j|~\�)�B������I�����G6�+�.@C}˻�������J4Q2(����V��-�)I����V���O�G^���`�"�_�%�F-b�[��\[%ț3�x�[��}��&��{�-�h4�a�aTk��Т�	�b��u�x�h}с�MP(v�K����E)!�i���q1�~�~h�r�5��d��@��/�]�xX�����.�%� ��ZB�ZYz�t�"��L���0eH�f�#?6���}���\�>đ��+F��d�U:N6��NX�	9�t�OŐ~M�J�x��wԾ ��aI}W&�$��]��K�y�9Г.ƫ��k�C����^w�,�M�!8P�	����g�B��V7�0b��!C�����&����)b=5`�U]���1�D�fb(�������-qd;�C���N�%�%��w�ɶ��f��Y�R�Њ��.]�1r�����!�#�F�7Dx�yy�4]�E�{��֣Α�N��*g�����F"��V��6�Q�q�� �V�j��˟,ē���H46��i�r��~k1d���oP=ۺ#�'c%I��En�<��	�.;�L4�G�+�.a�~�El�����9~�IυT��n=�l�{NCI5^޽��/�b���X��<�C�ZX�]a/�W�a~+^�Ulh�C�۽��_��ӝ���f ��ϔp�P��7&�kܥ_P����Q��)��w��YZ;���3"p����m�<gS��/�(�hc&jp҅��Px�ױx��w����>}Y��mmϧ3
�z1��E+A����^^�[?�`Խ�!��d~��<���ʦ�D���Sّ87�t�x[��҈5��=6�]�m�آ�^��G�E���Q̤I�;U��숏v('�A��`���g�A�*8E;��88¦�t7r�Gt�<mj	#=��f��q�́��!��z�~���Dd��C�f\��s�ɖ�����t�W5w�k`5s���{�/7c�hBQ�/m�Q����'|�t���X��^�L����{�ξ��ˑ��ζ|�;��l�.���]�`�$�:V-���$oɘ���iw]��x��A՝ENj��.fn�#g$9l��b�+��H�gE �-!ҳ��иP�m����'r��5f�#���389G�m��M;���ҫ��jP�Oy�o����'@���ݣk�M6p�Izzv|̴J�Ȯ/���R�boxDK���\����w<�֥<��%�!������va�`�ợC�a���ԭވh��b+&�4��ذ�f���G�hs�P���I����x�m�"�.}:'♭F�F�S�~֚є�ʆ��)j���뒥�ȕ5L]�}��R	4�}�xLyN�H1,+�(��v��5��[E���)r�'��L���_������|� ��pQH�n�X��6�)�S��S���)��~�1tU�� 1��q`W'P�/��v p~��?��Ir�txT� Qz��>�Ӏ o�0�)�CN�������yp0&�q�`���� �A7����y��$oc���Q]5��� x���o��(��}y? @���eW��4��|��D��A�7@���T���g�� ��EDE���3(�rR�u+6��!���������CX�1�aL뾠��f `s`��,Ӫ��M֗��h�@"#����s+(�z��Ϯkr+��Ű�e���=�N�l�p�t��I�(Q�,[�
8��kt�<��H��ܳ���wy��^��M��d���o�EPT������܃�*��y��S~�+ns����&�i�e�
�	��Н.?�Z����L�W�'�N[Wb����`��5�w����t!����@�a�خ�����V�ԥ���*�&�g�����C������1#�7�s�-��6K�%,U�?��YL�ͅ�ȧ�7��n�������-a��H�ƂQ��I��X������c(�mi9�c��J���'��,�yr&]��/<��:N����s����$�;o�b��ۿ|��ߓ���60p8D�F<1/2��X�3t�{	"t�`kX1�"y4�P�k?�1����ƝwJfw�.��8����^��l�l�)�\�)���X�+�����z��`q/�|����� ����Ѩ2��\��#��Xp�S�X��?�	%�6�]��E�)�*�'�t���.�g�T��j�	$B���Y�L�048h��H���y��ߤnE%} ~Чb6�!UᲚo�t�[vEW�ǂCc�sBT[��@R�������c�02�"��>z�8�Z�]Z�;XP���X�H�e��Z�4���6Y��U�ƱEͪ�X/mᰣ�f#Qc��Bh����=�Ǐ2��e쀾��%�x�u��3���P�֣��<)u�Xxza]0\��������0�g��d��X�.�g�A+Iu���G$��['镭v�X��H�#�7a�.Ì0-'�(4��,���4O0P�ɭdQ�������[�K6*d]��j򏭼�`);p8�&�ۣ�De�#f��A�p���¼�U�<�V���a���4z�~d���dz��b�v$B�����4��_��OIt����eW�G�mC��p`h��c}Z�u�4�4*�	{����2A5^�)f��N�ys�,�[�D�17�hqy� �x��H1�U�pq�I��R�%V��:	���e���Д]=�B����y���W��%Ld-坽�P?���)��PǦ?��xx�$k��5}�5ԏ4��5	��2w�>����2̏o�%�������Ǎ*���:<�iZv�=P�S���-���
p i�˳y
cg��B�V|GtBI��6Z�~���bU�7��_�K"���@T;��}��x�$�R�~IzEɢeż\����osc��v��ry���m�<���9�#��5�AǕ<z�$�����1*�=E76/v͢%�h/����_�4E��elG�K#W���m3�(��D&�X�;��zd
�f�<�0��O��}������9%N��rRѴhK;�B�(�f�7�n|*���׆[��+��	D^qYz-5�7P\�
i9E'=X�fM�i��U8�|rJiG�TI�j.���p�V^Ӕ�\�?6R.d3+#�i;P��F����r�Ԍ<����{v�T�%��o4֤�Ѥ�E����:�ӊ��A���!� �\~L'el�0�O��_�m��C���+��Lmn����6Z��:����W;j�Z�H�5�oI� �`��]���2���|�����Q���"��{�+�Z�����yލ�_.��*������Lc�w.}fd��<���
��e��m=��8�-Ӿ����j�� ���{=�ϓ��he_��2vQ��b��)`f�T+��]ptg�� �'��Wٶ��������L[C3�v��e���;4�6��3����I�U�� ��V�O�Y���d�4���=�
����t}=kZ��姡(&�i#5]u�F�vt�t�䨯���B�K���@�F�\�?��ߟj9f��8,Ț�:RIi��X���ҋ��=���i�%ʓ���8g�Z��LTW�����͊q�j�l��S53��Z�Eه��S&,w糅H�t�H)��<�՚����`k:�́ܬ��I�<u4�Z �������Z���cI���/�fw3yc<9��f�<q�}2=����)^(Q�PG����Yį����m�u�9E�I�XE�+U����h8,�On=�H����|`�x�"�|� ���[YSO��K֨&d--\'c�p�,c1�c�`��xƅ�	�ia���S(/�q��0��-��g����mm�9�[\��&7��<�8UW�[��ʢ3�Ӆ�7�aV��H��n~����~7UAl��*�-�.�R�#��|_����DFfx4Q;��d�.p�^�tV�P$x�����I�ʾ��X�W�~~��n�U!~�<��DZ��8:_x ��MˈI?<��n:8���yn�~��?� ���Y(�%�;<�ب�qH���[=1*�i�ef���Sl;�|;lz���S�Q�����y��pF��f�3�ǜ�	gh<�-y\/p,�(O2���C`�z���Ϊ N�B���o?{��Q�yGLZ8�s�(���h��\'?�`�D�U������Ɛ7-`$W�I��Pp��^�7�t�6����&�X"ʜ�{��w�+�z��e�R�cAS�5]��m(ԗ����O�-f��������6����pr( T=A��w��'�����i�jl�:�ȯXy��R5
�{�x_���T\�u6�x�"c֐�,��ޙONp:������%H�*�`@�m�	�By�Ro}�{0L�.V�U"I� �6,Jnp�񚑉J��������3��A�+w�ġJ��������Y����*K&�'���r�v������ܺ���c&c-����X
a��k�xY�!��,��+`�n��X|�~'	W�Ъ�19�`��d�]����z���3=WQ���i�ܩ�gc�B]���r8���չ_靷�Э#�ġs���,�C�<D���-�+IN�:Gl�Mԩw �w�X�i${a��;w�u�u�6�&�n�$��e��_Ͽ%�PlFЖr���#���Tղj��tY4Z�XDu����G����(��߸!aS��;�����%�9f�N��\',��a,t0�}�"�]�s�y��k�p6�Q��xX f�B�
�V��W;Ջ`}V_�i�U���s1��'��F��,x7��C�9Vl�uY�?\��@n����,B1[��$w�3�78�[5~c}Ф�N7�^�7n�m0u��l�~7r|ӄ-#�MSjy_���X�:S��j��b�d�gS�
�#E�A��ݣ��ui�u��#!���[����	�ɡ�fBO�n��<w�-�c�9w���ZH������T]as܅u�DVN�gѺOl���t疲L��ּ%[[���!o��SL�CkC�6Y�U���s�!N����DI(Oҭb� ���w�D�-Wΐ+׬=W�b@eb(���[�v�U��:N�#�J�m��hȆ2$���[�t� �$��<����۷�AH
=�;��Z�d"���<軕���ߤ�/#3�P���NIY��V��v;5�S�(�ؒ�ȩ�o�^��Yo��A5��Mm;�������aՑ;���3�R�A��+W��.z���,k��]T�Ij�W�d"�c�s9{8�_2T�-+�q�A���'%�g�u�� PK   
��TB��(�  /   images/31ebd35d-3137-4c9c-9389-844452b616c5.pngĺSs.\-۶m۶m�6W�d�v�b۶�'�m��ۧ�o8����Fu�ѣ�f���$<����
�����U  �B%95���_R2�ŹI
*r
���UjZJ*Jr

*j��ե�����bR���������IT4t"bbN�nV�N::�
rrRPjj�z�鉑��Qz�nj
�n\\<jZ���Yv�.��^,l|�>f�>Z
�v�Υ�ŕ��Қ&��ޕ����:�6xxxn���p�3�l�]L�}c3,,,5-]�PH����Y)�''K�Ɔ�<�:��G׻�R���FfZ�J:���[ۛ���F���v��L�u6V��v��u6W�Qpr�ZXٶuL�7T�`��T��z�9���D&t�)�jx���lIH˂���M-ז���7�F��&tT�<>>��GV�{w�&$h��m�����99=-N�,(�7�:�S=RR�[<0=�5��֡�;���**X����<0�����Ĉ�\O�&moΧ�Ϗ1MD$-&��y�)o�+������[�����DR񄞡��h�?Bε�ܑ��h��3�#蛷4�go�׭X�����,�s�-�}/E������wp9�ݦ�������������v['���1tz�+����������2��~����Y������T�L��)���wro�����X������jK��e`���=�Y�E�H�t�$dd���������������$�~�?�?@���6�4LH�}���$��K����=�����x��ckcm�{�ܺ%{γ˻K�>dWC���p{�ٞ{�8Ѩ��>:H>vo�3E V�l��=��4-NB^B�x�Ԟ��U���|�h������揝F��;��{�r��9=��ݍO!0��k-������\���ݽ\�y���|>���;yz�N}_��z�:z8��ڵ\~~����l�n���12`��`�.ƣ���sZV�8W/-��.�m����o�Mw){�8�GS�n��̧�V4�O�OG�W,i�=���p�l�?�00Q4����j�؟&�y�B�xě=a�ܶi���w�N�h͞y�jŅ;�u]��nbf��͹�8�~��ڰ����xT���;{�S�<�6V�B��ڝuP����ٸ���	��ݺ�t�hs�$�����h#./�X,��pe*�!��	x~Rו����>�]N	[H��P��%p=��7Gv��6?�^��0S��EW�
~���Kt?a�>�r[XB��h�{Y�fMsL�=����7EY 4aAZ�5�4L�wm4۴�4��Z�SMa��)�v�_���'�~bp����:v�I���2m8�ʴ�p�� ����������p��W�Rw*Ϯ ���C�����Q��i1���M�~=�Pu���ef�s���PK"P\�+��[r�7�HR�]�x�*�ϲ\�3+l,42��|�?wP�)Oj��:|���"�J�`��x1;%h��<��MX����,T�׸�{����4y0��7�ͣ�^�&�p䈥��=�- ���KC��'�b��}�s�^�K�tM�$;��'a]�/�o��bfI켾�A<�'��Z�T�|&ԠC�^.�A���E�>�T!ln�4R|6�l�P�K��B����M<�m�i���LB�ue��ȏnt)����cF�(W�(l�WZ����o#�F�ow�D#=�l�\�ŧ����c�{�8����Ň��{����u. y##���߫>^�X�SDʧ^���UN�˝�����دƞ"�)�[V&ZH��FM����tx%H�ے����������l!eAK����s��la��Z�,�g��%J'?�eg�����<闙*r���1z�65��-wK���8R��i1��X��Gf�)�M��c�V�b�k6��l��!��[���臨#xм�P��8k7�c!	��:q�y��q�]z��t�Pր��at�V��7���]"��uKW,EC�VQ�ݫ�h�{Q�ĥv����+%&�VKZT�b�,�Ƒ0b[d���y4�Q������C�q�3�"�?x0�ѕ�u�������n�N��c��?➢O��1��i?'\T�D*:/��,p;���6��Z��H�@YZĶQ3d}5�i'����mO�k
��6#w����{^�'�ͧ��`z��s����"������{�̮�=��뚡NP/E���h�٣��@��2 ��l\���aߑ�6�bNZl,�6�}���!��E����.	��)T`Y�F��o�O��gkY�K?�t�Q5Y�FUtxP|��;�G�}</&m�{�{�5���O9���M�> ����UϤ,QQNu4Ql�-���!�/����r^�Z�N&Z09�R���Ǝ�~�*����&ڍ=<�]�-o/�O_�4�Dy/!�J��"MAe�߲�`��n5~�-��沌Y��4{�,��xkc\�9�r�A�,ȶ;�M���Bh�3U�ɻ��!=0�n�r�v1��{���[�2�!x���nqGF���
�bti.�L����c��奏B�L}�+������*|���ҙT����п9�������6<Rݳ��C���[z�z�A/���x����0����^8��XY���_D���uzxԧ7��!�H���/T�?K&�,�҈�al�1< g�U8
5��,��R�n��/]�;���o}� v@��p�������l�IzR�����j3M\�b�4D3�P���N�2Dh�%�$l�Nx�p�����h�q��:�@�*��y�⭑Ls�a��/PN�p.ِ� �jvbDŜ��@A�/<�"E� L+��C��Z���~,q1���CȌ��4�s����e��J�e�O�!f��)sgAC���Cr.�9ë��!sP8쩰2��mè�-������o��[F�	&�f*�i����y4��z��=N���[¥�We=s^9�I
+���jP
{
�&�.��d�� ���_�7XD�������X������j�'�;/>�Ff�ؓ�)s:�_�!e��C���J�r֢������cӂ`� ��Wa:Yu��S�]B�!�� Gc��3���͜�(D	��q��ݟG��)]`�w3�r&�S9�ԏ~�h�,;�)��슒|c���NĽEQ�r6/�R�"�Mæ'�+�7�@U���~��o̥p��`�����5��~y�W�ˤ����6w�h@*P[����w�R���8�d�
�S:���L�� V' �d��t��s�
㢧����
&��n��+[��K!5�������+����}���Dۮ"�t���O�)�	6��9�/���	��ə5k�����q"����q-@���Ո��d�G�⅀ �Wb����m}�-��@ �!��=��h�~v��  �_g��� ���jS��O��l8_9����#%��7G��v��P���]�+'d�[��^6],�i'�)�|N��$��^7f--Q%��8�����>-��vS7�];�g��2[��:�!p�m[�w��}�9X+�	ސn�! ������A�9�l=Ba����4��A��� gP�o5�;��S;�a�0$�n$|��ꛯ�+�/NXdGN\d���V��,F�x"Љ�vm�S�	=��>댯[�}�"� A�WדW?U�Clk���]�}[�l�aE�����0�ƄW�����7�I��k��G\����T�&sJCǤ���a�W�#�L���N������)��-��q�$@�ek->`=�\���K=`��v*)GU��2s�X��Z�eҲ�zq�-	�������MZ���4$W��'}������vP}�C��$zh������Ee��1ET���5��>��YE8��lr�ƹ���
��4�:�V�D��s.�Ռ*l�����s�?��K���	p���ӗ���,G䵞\_�?L����=p��B7������$�HǬr��az�O\�7����>��#ض� �T �eO!G҄q_����M�.Ӫ_��tR��Q'~Āv��Xm�b���S���}z�g��.�>�il���:Q�s�|(��h�ټ�)��IrNg"�����lBA�Dj����aXC�_`g�<�QHo����6���G��1��N׽L�Qn��+FY�w�Ø�74CY&h*�B��4\�)#!%���j)�l�Ķ���;e���o��6`�20��?S�-��}��y��,�1"p�ߟ�r8N��1�x�	��OPn��٦S~N�D�
�.��?�k�?ٳNc����8�������<�"��><.�	d��J?�����d��?�������N��GXҽ]U�)7�"�˸9�P�F�ք��?�����]rc���wcB�v�u�(f.���\?�?�>�X�Y2�$�y�u��UX��I�<�R���r���F}iP7��~�l2�`�-�T�v�.<��&�`��S�9�hi����TfO�\t霨�q��)k��M�����I(�w�������i�H����{�$T �C�]MP�2r��|�	>�z��=V=vh���8ӫ�������";ޥ�t|���̎s� p�&�jr�ͤ̚��FƶN]/�4鱐m-yp��۷�6p��2̝6q�����pte	�5mxq�%�5�������'ԍ�f���bH���1:<�����Y�~��ukm`ƌ�w��]�)ꦟ�U����i�*;>x�v�yp�ɕs�Y,���n��*L�6�7�������=���'����������4���B��&%i��cԓ�d�}\jRj�l��yW�x�Π�݄fK���P3GL9�UW/^8���F��G���]-$����^y��c�R ��Ψ�/����9+WAҔQ�~��N�I�:~�2�V�Ѭ�	�`71�����ޙ�����ur��е6�)�6۷�����d�w��.�]l�(����
�p��]nq�'Ͳ�o�!���bK���9pK�V#�+��}��`{�jn�,Q;	n-��p�����G�W���ȓ�^-��R�BpGC�ƌ���
����A�<{"�֦��
�^�������d�2M+�?��J:فB��W���j
uF�ˇ�J
i�/��_w��,1q*s'�EZ��3�?s;ݣId�9dK��RZ�h+�TN%�ZH��KƐ������|!a�����3y`��=���s������f��Q>�bb��5o�_�셱��%���k�d����<��������3��u���߹� KCKc}��K��ޭ�b�[qC�׋[���g��R3iV��=}�~��\�)z�cZ���5Z���IT7���_#�<�>���N1s�ό\CJ&�N�SY��L:m�H3��]G=�Y�Z�D����M��s5̭u����8�ܥ�#s�.<�07��	�q��bk�9��A��_N^�bv�Wk���f8=�����"��*��@����r��4+���m�s��OkO�3����ߏ!�k�k�*�-iIb��畟U�7>��$�Ů(�hM��^sH@E��͝ݯ����<	ؤ��*Ԗ�	#͈�Z��6\�ɧ�ݔ��$�O!�%WO!�HCڸ��%G53�lL�I�E snمU���"^�>��@��;�dm��� F����}C/������oe8b�Sݐם�)b�Q[�׫��AqA�U����R����c�g��E�7�%W����f��A-Ek�)R���P�����g�i�	��Y� �g��N{��=�
�$��Yψ���F8�!LǏ����	��G�'�.����*�����P����8-2��=��@S�*�����r������t���p���+$u�`71�<@�x�C�cCeU6�F��TG�ݏ�/�R���'��r
�;>*~3o��T���t�B��W��ǀ�5��a�qQ���W�~��2�����6�$�d���y��"��a&�܀�$�v��*:AÂF�H^� F���4dl�][�{C���g��8�m.+k>����p;��2��_7�=Lqa��!,�*/R�26F�9k�Č��5����c9u氼����w�Y'�!֯�I~����,��
7'w]%8�L�2��#p�d�9�<T�����ܙ}�ڏM�p�Z��U��{��n=wn_�n�)Uª�e�V́�&J)��m2��E� ,D����s
����[�K���C�Ӻ�M���zcq�$ȀQ���&�1=����~�A���P����>��Ѱq�|��)�A���h�Ī��OYJ��o~����b��	�r��<2ٝ��$�瞠h�¨�B�`w*�qF䜰�9�&3$%��iɛ�t.��y?Cx(
��/
�_!�0*��o�|�4~f��WJ�=�%�||��@U�����)Ә�J�R�yN�ks0@E6V&J�Ӊ�粡b!�I��?�hg����`�ѴY@_��� ٸ���ˁT�=8����ׁ�N�����Q�.l�,j�'�Ƅ�x���n�J.%����F��z�#V���i���S����.)M�G+�����?�Zsa�|_��'�I0FL�O�Ǩ�V�m��J��z�'�%ݨ�ȇn������R�ꮺ
�z::6N;g{��F��0�S��N��SB�^�ɊH:��d����k�c�g*a��C�O`d��ϐG���5VW��O ᗉ��m�?�A����'�V8B�_�����oX��ὔ�a�q�X����L��F\�H��HES���{����ش�8*�]���>`ށp�B�tT�t��M�����V��#�AĒ/���v���h�#o���J^�?E웣�F/�B��'|�Lo#����<�l�*[͡�� -�l��i��<զ��B�8':�b���w����n�OϢ�7���yh�> �5���$����J�E�����������O������:����5���dWX�x��b�:P0���0r�_c}���>f�����2��-C����Y\K��j��ˡ=��o{6��]���V�g�u}^�F���Ҫ899�~yM�L۔ܓ��À'�40i���"ӳsaф!�2f�rz����,&�U8M���ᑌ����1aG�u�]Ù̆���ϐ�"m��6�.��=$Y��gzU�:6HRb�������ɉ��G��$�/�w�м$�<�u�����y�c�c���s�������;�L�����e�������nO�	wn^w�?D�%CN��kz�>Su����r�0�g�/GBζ{��[���*̵~]��ɻ��lN�3�_p�;�p�9�t��v;*),O�,W�5�����?�޺k���X��7I���ʕ�t������.Ŷ��1�}�Ko�S��*�������������i&.������y[4��+QzQ* ��>�p�G�I�_%�p)�BH�!����T;��[ذ���흫��n=+@�5��ǽ���f��9y̹��9.���ٞ{[��vbI�\m�&݈�b�8E�u�fi�jR
3-��.9�������q�џ���ҲB��J�]�xLa�e�z(;��Hs�cƧ��]��%h�칮�>؁���^�l;
�k���6��[��e��z����(ʑH7���P"�P�w*��6
U!��ST�Gg�Xy%��d�ٜ��a��	�����p����
	~�~w�*���LTyc�,�_�� ��=��'�D�b�o���x�^�]y��9��đk���Z^�E�FnE���o	�����0��2e#Opć��`��g8��u���L��O����pY�FR��_��3�����+�[p�n�N��	<�\��]�� �<�z6�{&��J9���Ə��(Z��K ؛d�tr�2~��N�q��!�a�&�:Qg�Q��.�S�i����e�7�Xb��V��ElzP�#���W�2w�t��s&9����a»�����|.���X���1�*���d/�ES]q8u�;�6Qf�[�aW"�Z��5�;��2�
��&?-�S�2\n��s@��z��@ �㐽�:�.��E���w��+��_P�ZUDz�+0#6�rߗ�X���r`Bl�M���˜g��X��c�Xg�ځ��^[D2 !S���b��`E�E�".8��u��菼����͜�U���W0�:�1�;�i��/�<?|��N��j_�\��*�[���.Z����1���n�ߧ���:���n�pp�/�X�T���M�$u�sgKx:`��w�Xb�?c+�]�����@�g���g]\(U@#Շ^���zi���V�\v
X�(�R���7wB����jI���lxו�����4h�����Xiˏ��SG�-���r��h�^�f���������7�|vu��yk��'���DK-�s�����hQV���WetD�j�i�e���گ�
T��ցvl9���pG/�n�U�*�V�RZ螴Ӗ�5��: l��|�Uc�e��&G)�G�s���y�LE�����4=v\u��&į����n�r�<�Q��&���  ���qb=cA&*)$̇M�Q�����gµ*�}|ݽ(��Gj$��r1`����G}=$?>v^*Jj�
����t"'ͮ��r�U�pM�82s�>G�l-:��|U��q��ڲ0G���ҜU�.�S��8D���[
��Ds �m����lC>�>��z	�����ޑ��{ZP����p{oLea�ה��sus���tu/`|�Ǆ�?f�G}j��U���1��3|�4NO�L/�֍'�P�&>U����l!_ʻ>���ǎ�w���w�r{���wۺ�\5���{h�~�b�7U��k[ �0B�c�pN����E�-�,4.�=��U��GP
��\r�j��X��n���g-U�]^,��BD]��peʄp��3���4")%�c�zȔ��O����	������Hpס�|}�9�T�w��(=�:�A�:
�leL�_�'d����	��D��3�W�:D|J�����s.�������OY�߯�W�7]*�4��-h+��'���������W�Y���T�]���<�z��~����2��ǿ�`J��E�J�Oͣ�֝`�^���KQ|��.T��u`�\����:�\�T�r�:`��N�9�^ևA:�dmE`�c@}�0�(��ip�U`
��0�r}��߃�YR`8���Bu��|>��n�[ؾY&�_�� �Ze-��?m��kW�Cb�0<"�$ᅒ�a�4T�O�oF�-¬#���r�U�ꂇ|��K�ߞ�6%�?��@���<3��N�ދ+�pg��.�h�+����	��Z�O���w��H����{�2782(g�v��M8���+�^�\2��ũV��'���
��F�O�j�J���;���.�	��﬛��_���q��U��ݯ������Y����� B3�h�y�'�o �<gz3�I�4ڍ�������Z��L̶J�����^���5ӂ̝vn� ��E�̮����i<��v�l�jT��6�Xg, �B�I;i\��� y�t[�W��@A�N;3�C�ú���(��4ס;K�x��`!:���ܪ��sT�l�=�
��qI����K�����5�5�Yu��=<损����O(w������K��E:���]]�MO��c}q�U-l�J��勂����`3a��S��C#K�X��W(�3��s������.�䄶Y�wfVrmF^���ڮ��~�(;p������hJ��]�`_��� 2Z�4w���e�F�8;�5ĥ�M:l`�	�f�_�eu�uz>zs��܊h1J��J`����3|��`	(�� 盋���������󯣡���������-�!����n}2] ��b��OO�(w�i,�.H��y�rڔH�*�/�K�F`��K�����ޝ�b��+��Gn�F����� }��/��Eӹ�D�k��O�v}��	@�����8h����La,��|�D�~��O�A�{����w'l���k��UZ^���뗖 �<�m������vm �A�a;�[�ɣS8�*�������\��gO5��jk�a$J��ճP]��d��V]NGx@P����ԓ�rŘYI�Cʽ�����oq�!�p���Oϴ~]sA]��F4Q����&�ɤ��+4��g���b������*f��u.~�u\Vƃ�[���nZ����lH��hd.k��RK1�U];�v�����߻{do��c��������2��R���|�|���6��<am�\����^�/��S���L���!��Ã	�*�� ���^��T�5-<��;i=�CUL�Q���<z<�����RӉ\��Q�v��c%3"Z�G�S������<���Bc���t);����B��½���z"�sc��9��a�����x�+�k����FQ��J�97���xjH��ӥ�yGb�K�?��R\r��f����������f-�$�N�Iv�A8{�|��7x�Ԧ_��ܱ�q�-Kp�t��ӑ�Cnn���N�V�z��u0�5elB�=�*���9��P1o�U���r1)�)[�A�.@�Ê���`�p�P*�^؂�%�;@�;��+��l��w���
�h�.��L>�eXc�W��"�ιE�%&�7V;S���S;���£�c�	�[���!S�~��?Oπ�&�( �m����Gbn�|a;�-)�����x�'�$�\#2�j=x�m�����'��l����^�ge���RW��S`� ƙj�t��� W��+�܀�ߧ!/�'.+Y+��0VK��>�����~�Ev��f	6z�����xy�.� ��<L+��
��^��J:�+X�I�Wp�۬ǡ��1�}z�޴	�5{������\�lO�.�L���R�)����E�w����.���@	G�.�E���_�r��y�v�tĸ��*u�v��x[��y�n���TCGu��� �B�����|�M\�^�ɢ�ԀF��)�blr�4h}jJ�����-R7�n��DN���gQ`B�?G�,<��a��
:<��m��F��8
���(��A��=*��(HN�Ȥ@��؄ά:x�G�a�k�g�a�
�Zhc|��!�J�����$�(u�C��H5��A�iΓ�0������vK1�|xL��W� ��
24}�_�{J���F��,hy��k���ɏG�р9�}�*�DǴ�4�TԡR�}���As)T��.˚e��T,�))���E6�3��(d�rL?�.s(�Gm ��������:���o��w_��jX�����+�T�	$�U(x�I:���r�;��y[�Ru�%HZ��r��j���;�S�#���Z�'�� �D�Yx���(ϸ���́�I�w�4�6aǚ��_���5J/��F��Vv$NE�����?\�F��ݧ����x�*J�k�
u�Y)��гl{�t���{^�TZV�rF��l���H����MhC,xY�m�:�G��d�$2@�AKAV���XZ����`���S��f��w�j\.�a�T��24A ��SPwJ���
���[Z����$�@'n�c��Q@�Y�TF����&'cX	�GS*K��sa��'g��KЪ��q?��2[v��qL��G9�Q}�G�LV� B���I��2�A@��mVP!���8J�@����\��=����F$F����J�cz�-G'��j���H%LД�S?�K�-6�d:X�`�
Ȥ�G:�,�����":�ϴ��2��t�v|ᗬ�X��˧��LE����5�ͣl����JN���K����GJ=sn�Q�K,����U��Z}ז�����[�$�A�S��~���)�|aJ�+m�,4>LJ�v���<M,�E�[�!Y�����0����,�Y7����F���s?��1��A��|J��~�E�:�� �X�	W����Gq�w \�pJyX|�Iײ�����x��U��@RI�xU��+^����4B_�r�b��8_G�a��O$[L�_�L�˞D]s����MXV������\q1�m�u�~�J�[�u~�il�7�#��A���u5E�u�m��N���O�q-��~��M��ڙ�TWM-ʐ�r@n͂M��N��w�Z���	T�Cs#�q�Y%�)����9�!i����RS��$��y+3�).c٧��������b!�����ס�׵���9�h'���^��aK*T��VꈘE�2@�ٖ}��1ȁvJ�Z]B4ߛ�C\ܢ�$<����ȮɗG˒�À�@^TK����Z��
��:��nUXє���ZW�ͽ�d
��,�H�nʨ�D�g�7��56a��DQ�������r�l�����L�VI��a�^~c��uN�n�K��Rp7����hλ�����ߝN0�x�1������W�����DRī�E2�ސ�B#���IG4e�?y�x"�%��R�;�0qU{��`n��Q_^�1�rR��w�Ձr'A�<\Y�W;ҍ<*�o���T�Vs�5�sO�F�y6	���sX���{g�#n��>a��Wq��n~΂�}��Yy��:	�9[���R��%�����S��m���i�Q6x�qw!5���M�Y��Dٰ]�Dq7�7VX��Hܴ�$��Dvk�UQ}��|
�S��� uI9e�_J�.����qV�Uy���k��_,�=pd��H�W2��ɛ-�S�O8@�r3e�%2��9�h�`�9Z.����Әܳ�H2W=Z���N��8:�$Sj�7#m��ʥR��ؐ�kw[��ضd�{���Oگ��q���C�|1���s��Fw�%@�x���(�x�"��p���Ǜد�[�¤����"6Ũy';/XP�Z��jY���
��ʝP�1�x�eE�אJ�ƮK6`�p�:�<����sr����z����0�����7�y顺���
H�	�e*��ڰ����t���2���2���O_{�?����kU��eT��~��+�y��TR�j�><7}h�궫o��(�����.ê�SK���&�	�Pbkk����)!���A6��6�:ΣE�ދ�f�7<D�����nA�D�j�;f8��(� ��2p��m��χN�*���;�e?�t�% ��-���L��bF�\r0���@/G��]���B���"r��������' ��3��x�4�>��f��I���l>�GB���ֲQ��6ʴ�tZ�]�2�MM�?�	��22���ϥ?�z����t�����M��OMM�_�L���D�s�(�#�?�so��U��m����:�~��T�?�|^�|��zz���\�慳��UؖS*�X;�ZtqW�ɐ����+~=,��?������z*y�+�g�l6A
����6�9De���[9g��6�\R,ǳ<|̝�B8R�(�3��L�^���?�
�(_��9`�������(0`��׋���S�A5��w��	����}�\��Lb���
��s󏢔6p�7X���պG�t�v#����?�� m����V�*;����ݓTWӓ�ŝ��e`�����e�lp�a������ʿ�a�w�������u]�V��m�^�_:L�c�+�Wzɑj�h��p ���a2�v��s|ӉDP9�8���Q� �?k�}΋=�4ϲ�L�����Qo�c^'x}��2@n� � �X�<е�>*�j�M2Lbt�k��M��������� �a�#�6i�f�3�v��Yqr*)��S�<�A/7��%��CK>���/>\�Q|�Vӭe �V>�Mr��~tQ�ݱ��p��q�(Tu��<w���=6���t�/����2�O6�5��O4pC��@����7�س������� s��Coz1�ӶB��X��Pp�9�,3!�8�wb�ԍ�ky�(�2��CPoA� ���Ϛ�\��1�I��[����+g�F����㩬B���/�f@�QK���mMͧ��W�д ���#-����(ͱ�U�h�8�@�j�`W�m�Z�ak�m�#�u���;�VR��2��W�Bǣ<^����'�v�O�އ�%�r%���S�c<4k��	.c�6"l���弙��-Q����D��'�ñ��r��ɣP�*�3��^�-�f�1!��P����|��ORS�p^�ߍ��ӡ9� �|�Ҕ�$9AΘ�y��ϣ�-����l�/�$�>�G"D����p��$�oQ���q�E\V��0
Oo/[��k�J��`�%e�����3>ff�t!-���+\�$Mt��Ņ���n˨��p��˟������5���bV�(����p΋UIݱr<�u��,�}���n>�����ov=SzNo�_����8���	�95�v��e����Lf�ʝ���!��GkS���!��4�b:H)9�Q{�
��ND)� z��~c|�e��d�w�%w#e2�/��S�]9�"��f�%�g��m�0��-�{�CB������`A�Y�v_ySU�������P���W�Ѩ|�"ɒ!:�����n]ɜ���3��7F�Z����6��N��Հnd���ϰα�\τ�P�ظ(�G��w���Tדm���B��~3�Ff���އ�N\��	k��T����{������w���`��Ѹ�^D��.��	v��z��ˀ��9E�u�����9+W_��fWc��Z���>?�]�8��u��)t"/��5��}x��G����+�<ʤ u�qU�{X�(���x��.1��KlS�}O�J��+6����b����)�m=�ŗ�!�̓�B�s|��8/��2Rq�s��5�1_�����/�C����"��W&V���a �|�����b�"*,�c�y̧�'kV
�^���V�aU��#�8���Ch̅�Ut��j�Ì:�@�eU4G~"����ʈ"���˵w��s�P������b���S�(U���Zi���KX�fnC�+����=��m ��V�ɹ���F�ܷ���\G3�TՁtF��*h ������B�i�M/��ͱ�/��p&]�Ώ���	�*j<Yђ���n��qq^>����d8�G��l+[�y��O�+���~^I�~IJd������k��ձ��S ��IP�:��а�/��4w��3����m�m��"�8���%������V4�Jܓl��d����m����=Q��"�G
�5*1��oJ�\���ؖ�l�)�ju	"5�6��E�&���c�o�4v���!���E��0��JciC������5�j?sf?�ԛ�W����Y��|"�bč��=S�Q`�C�U�bʣ�G���}g��ܮ!�`A���o��rQ��L��ܑ������2�*�R��4E�&�?ɼ��N�<���[2@B�뱪�ݰ,�j����WJ�b>�4��p3
����F���+�07@��>���_YCmS@bWZ�/��6�8\�;^B�{���7Hi�.[bH�U�#<�#�j�U��d *����*&�l����v�Y��r��j�� IFJ~]�����ܗ:�_bݓW�9y��XJ|�G3J�ZC<'����}J�\��R�$&��Y)�lTv�Qh9�6�8��yl�Y:2#� )���Sɘ����e�a�Fʈ���L%VS�MJ�p�-�I�$���PR�<|�$J8�­e܇���q}�������*�[3����11��։��*��Qt�+� ������'��z�M�����6�D�"�-P>3ܛ�1��hv��Z�.Ô�j���f�@s8ꢛj��3�������O��ۏ4wS*e2Oƛ�/�ls�O2{�Ƿ/�B@� ����P5�i��r��{1hl�y}0�V�ٲ@�,M��r����Ԉ��ҫO��HLn*<�6���±���$;<������]ZҺ������K(`����Ǔ4Fh��\\����6Kz������	�ۨ!t{��Q1�9����v��z�tQ�0Y�JP9q�(���R�ˣ:i��I�4��P�m߾߆��MW��)��O@W_���v(����w��
?��<P��9�ke�Χ��w�"�~?��g2Z�Ի�v��M�zW�Ns�?(�C�{%��	�$�����\F���B
k��*��D��%�
�kT���'�9��wx�6��=��ُ��+Wb��p�k���;�US���i4Y�-��5���=���S,����{ay97���ηj�
��;�R+z��\詺!p㴐y�o�1	_�r�I�Kmv���V�����D@��5�;�&�"�;4�e�F�:� �>ϫ����t��?ǂ�i��+�;�����l�{G���I�Y����XP�χG�{��5��8�ʻ�K0z��<_�t_.��	�r o�eHv� �9��P�G�r��T�8�Z�Q�J����ݍ���0�/Fi�� �b=��P�2lcQ�ℙާB6rV���7U?�裀���eC�+P� r�/��؊�zҥ��6%}�΀�����o1����θ��z ��yơ��UυF�,<̳Y�N���	O�	l�c����ҽ_�͠`�    IDATgO��}� ��T@��h��Y �L!\Ƕm�v�F�J���]�����oNΒ9`*U��ד���g�jJ�Z�\D��?��k��o�ˀ88�j�ޙ���/��	th��.fR��Y9�Vv��^�����O?/~������H��	���ӭ��^���$�u��yo�����Yҁ��@�
��5U&�V �n{��G�m��
��*N`������m�=��������07�ma�A宪�=�'�����A�z������e�������E�BL�,y)\�:��1�{��vǅ���G�v�ٞ����F
��>��;I��}^-b_�۬�����?^��st�L����V�\}{Z��/�
����_�.�k%�ȋ�U��^iT�5t#+4M+-��X����ƒ�b��q�k�oa)���b��/7���.����� d���688���I���
��
�*����R�''GI��!#7�cJ�:���
x۱�ٰv:�<�ڌ��0���*0
u!����ԝ})#f�I����E| �޷�#ԣ rlJÂ}�����8�&��� um�w�Ǳ���3��ڽ����8��P����^�̥;<7��2A,��_��/ww7��׀�2A�^F}uu.ݗJ:zq�W���\���ӫ9'�Z^�Y�q���=+��7��ӭ�#�G��*RƘ_m^Y�ң����;�9�Y�_�g�J��i��/���`U?2����wώ��/9c2#��j�@�p�Ϭ�~Ƕ#յl��h��+ggIwzt?R�y#*cN�<��s�ϫ�D�/�0�x6���FS��p�~���$��]A�����o��M�Ν���{��qP{.������������4� fO�{��:��p���o[�d�2�}Y�yJ���{�bN�xL>�IK0G��s�o���Ӥ�'�/֣=4�9Ќ�4�eg�9P$�Zz�pL����&=��יe������}���I F�Wҩ�G���O����LL��9���kn̼�,��nǮ n��N޷���wΘ ��v` ���aN�@�^��dٛ��a2½ϐ�#�+â;EE&�t���,���:�� Ň4}{�.�%��ïH�̫���m��~uy
�N�Y3�k-K�Z/���ps�����r��^�p_�l_���������?׊{����7dh�͐�}�jS�$�0�,¸�zL�Wy�lR1�8��3����ϳ9����s��u�ȴT�V��&�f��'�� �!�a�����b[�1-�G߿atve>�	�{2`![u�s0o�CUVɏ�����p8��@��aj�`z�� �}Q^��0.��H�\���Z2웢[�qT�	�r�z��G�Y�'b���d6���b�1͈�ݧ�f���l̈�U`�A����Y������4�i�g��o��<_'�ύ;�lˢ���/O.��4���y�,gM+?Ow7 �Y��l.��X�t]6����ݭ���0�d䲕P\_T)|�t��LWm��6K�~gx;}�#��0�6�cEUT�-p����'̓�(��d���G��:˲��AĊi���<�:h�I2M��-��E��ov������LA6*��,��}�=o�T,ј��^:8:����Otc �6�z`������Q^�N��,j���������ˢ�N�^=1�r����/7w77��- ���{M��,���;�֊EN�����RI2����^�hT�^]H��zL�7vX\��ᚱ����k0z���Kz��V2���~�x6�8>\��Cj.H�Yy0����c��Y�������M�%q�	�ΰ9��%г�����I��0&l��ѝʂ��>4�P�6�z���V�؟㿡t�x�����^%+.A�n3�=�����^�W��8�~M�&���8�m:�8�y��F�载���d]���ʻÓ��/��|N��3�������<|{�^^m�B�/�'v�������^�u��^]����-]Ҳ�}�s]VuM\͠=�9=3�*b���B�J=>�H:��� �V]Q�빮?N&�c�j{�F���x�D�| �q�1�M�]�Rp�C�&Ni��S�}	��]&���i�V3?{�y�ٟ����Du[��s�s�7��� �޷��^6��jYAo��uu�,m��bf^ゞﻞ�/S�閥8��Nܯ��;�?�#�M�
K�J��XVo�'�7S\!�3&�Q7_3w�'8�
,��98(�8���%�����ж#B���q���]�n�\��O���<���ˤ��ڝ��B~�������Gj���V�� .������ӓ���D:8]7�l&=�����y��5� ��G�=�����{1ݘ�7o<��^���Y#�8�\=WzR����l�Ç*�*jV=����g�������9K��V�s�ޔ�}�.�.].�ک ��-�2��37� ��gCsg��������Hk4t�P��K
�";�u=�ޜ��i����Q���q��:�s�2�^u��[�]K����t�m��O����)��
;ZXwo�����/��vߦvo�<Ma1irɗٽ��D_2t�`7��Zq�!����?4��̾�f�=2z�arwXZ[�(ݏ߲a�22�ؑ��x�!t��خk;��WU��-��L(��/&�'��.p|>z帖sx�y�=�J��.�Wf>K�UO�<r�$�Ĺ^���@W \�UB��TG�>��U^N���=��z�i�xѠ[�e���mwϋ@r�I�B�^�U7�a�]*ft��eCֵ�u&�'U��b+Ou�^XY��r{y��O�?���.�qe�[����Ͽ|<�}����:e�!er�:�q��/Vnp�΀>{�٣����)����ª;��%.4N�S�R��~�n��
�q6p��{�HN;�~����D*��d���2zќ�qcKXj>koVΙW�B*w'
E�J/춁K�#��ٸ��)��$Gӣ��I���I˒�uOd�'���cśT
,b��f��%�_��<�B�q�����սZ��u��3P��*=�>;�_#��y�y�P8�r�����w׬��H��$�����G/����%}NN/�5�ˍ�`�,�Fi��3�Ϟ�dt ]��u��ޯ<[�%v�%I�J�T.�IF�#O�V,��d���爐KFǇaO�(�m _�T�h��z"<z�[�u�m��q0acI :w�*���MϦglZ�O|���?�����Qo4��8��5��Ȥ�-�u��DU=r��?'��� v�q����g�]��;�ۘu��6���f����3��L� ��xS�.���~�������-1i���{�:�;<��&K��f89�����G��������g�=>��fƔ$�,�+;[5H���PԸq�0���՞�/�r�zm��SC��e9���x���C�� ����v�W齳�x����(�$��@r����h�mE���Ʉ�t�j}qw���x���~P돺�U��Q���qz����~�L�	#Ǎ�.<�oD!��dx����#;���0�{|��mJuC9Hw�����=�<��,��"��ї��>Z{�W('�lI����I	�H�?��-k6S[?	F׸}Y�g�}��/З䆩�fI�x\yT{��Vz`�h��r��g���%ͻ5ױ\�?�t�*� N��p�T�U:x�з6~����N�-�{�Scx�A��"x�m>�)�dq��s�c�FL�
�L�� ��.V�27޼�=����ˆ������
G���?����'� s�0�C�T�� �C�(w�F�����_�m'��2/���rkq��:bZ������[(�<�{��Xh�i�?�_���>y���`�l_��1Ŋ�e����zUK�iuY�f�>{�������r:�5�͝Ǐ*��b�y�[�Y��17�艁N�
�F6�4��@�I1��t�Yv���iU	D`F$�R�})���w��\��E��F3W-j�'�|2���n�U���V9�
a�Ÿ�Ĥ]V�T�Gߺ��x�:,������_x�����ǝw��Ї�#��(
� �}���pjd��a�sƃ���//����m-��V��,����c�������3���p�YyOf����d꒱ �2\�Z}�Oc�@3�}���o��'�k�n4R�������d�,��{��Ī{8�����fp�f��^|�я����A�����EAU�Mo�&�m(�b��ܭU�ģ	��(�"�y��!<�7a�y{0𪍗�9Sy ���z��R|R9v���{����cFan���'͹Nd;`�a��:�g`v'�9�S7��\�IbL-� L�hj�&��B�s�k�Тr��<�=����"3S(��¥?��~yyb@�S"Hs�.�8J/��+����,��)��g@�=�t�nBL.�;����k���T�L�@�Bi�{uwq�3��@g��;m����,�'��>��J`���Z��9]'��#���������܌�d�MY ಮ���;�Yu����(��p�8Wl���p�I��,��|�}C��
l��]W�tU���+'�g��u/�!�J+�"�I���	FO�s�����o��y1P��^W���|���5,�^k���6�������i]����Ε�l��Ƶ���+�5&qH���4)���D[J���@�"ѦH�vi�j���q����}�d����93g�`���{��b}��?��Ba������|���[^�;X�?Jy]2N����g���1fsF�J�N�rU�+Ii}�l=����$��6�"l3 �L��=��aLUul�tC
�(5�����q�T/!l.��)�:�	D6����+tYD��I�3^k�z(�Gh���1b�	��0G'�X�eϸ�a�17�L�.�q�o�>�dڭ�p������v����'ϧ�i]"�A���8��(�ӫ�j�bq���/��з����_Ig�HTݿ�^?CF�d=#R^�@0�r���r��`��������N2���g��鵂�Ɇ���$�khPgKh����/Z��Q�v���1E���6��Z�i���P�ڡ���IQ��c'�w�*Z�BV�@��(�/F���3�k] D�ѡ�7�dܩn����ư�#���{��t��,��]�����鿰�rb��.|fb�V����>:���+(H�xw� Z;����(��&��.t�6���ej%E�[do�"�d? �����_�!���ӭ�I/���/PF�z{|�Z��5����̻Y��3o��l&oԤ��$�'�>}�JНp���}��wV�����V���GpM'h��ئ�6<�V�����u� ���ט�4���&�k��|�5/�R��	�cC�B\��HE�n8j�ǽJ?���{��K��u �YO�ʖh��N����	l�q�)Cϣh�i�`��(;<�.`��q&���a���p�Y?�ZV��	sS��9�>Ga<�W̳4��^���n1��u�b�Fg?�9T�o߼V�� ��dLYMf�r���I�O��V�K�Q�,�PxX���ӽ2o$�r2�f��1v�G�ݡ������C�<p�w�TK}�����l.�bT��Ef��R����<��d+[�@���!��iƁJ�������8��Q�o�<xN���(��v�ʸ�}�f����1Z�*�L)�w?��� ���c:���1�A�3N:p�"h����b�eЧ�^���1����uG�=m�-�rf�Al�(:�Y0�zɿl��O�	�w6�ܼF՝]`�?����t�$,�Թ�db�p�$�'�9���!%��bme�8�Z2��3�,�55_O�?�X�F��I'r����x��G�葩�L�pe�X�	�7��~�1U�O���d\��=tT�ĵ@_L�h?�kw�Q���,�&�m�*}G�����r=~C���g�f�'1���+낟�t����i���{��	�HJdӇ�K!����e�o��`]7f_��:����R$�>������K���n�~{{tt��~���̱A$����^��z���(zF�u���k��we�n�j.7	�ɹo�^��a�ז{+�X�`T�'ܐ���#wv�\5].�ۈpdX��1'FT{x�P����1��&1_^4Qh�%P���5r��Q����G'C��;<~ѭA�}gHq�IZ�s'Rc�`��f�������U�?9'��J�1�����Y8�z'������ibAc�߇�6���9���A��4��@	Z�Gкo�e�{�C�������Ot������FZ�{A'��������;��,gVc�K�Fy^Ҵ�I�O�}B��V��z�Ж^�!�8`�U^�&fr�X������0vm�T!?����v1F���L���n {W%TB��G�j�[�.�;�d��+��,��"&���ǫ�myع�ݱ�+�v��Svy��G��Ó�~U��.#���lV�����k��� D���qv�k���`J��	�N�}:t��C7�OzP�Uޖ�"2����׽�m��;�0-�[\���5���}:O�7?=�{��`�.�g�k%��K"�^�����`������&�>9�y�>�4����ҋޫ��do�jM�S�U�$9k��ŵ��)�Uձc��N�9W �����a��0�u3P�J��D�p�q�#q��F�D�K����z8�~SS�m���c�����T�>?A�]+L��aB��5����@,b����>:�O-�m"����M2�)�Ch�	��۽>�d���PB̎����=�'X#fuY�em��Wo�_7y���~-�4��<~B9|kk�A/Xͼ�������5Ү����7�^S�<::\`��l��7)��t��M}r�7�KZ�041K}ck ��祬 �1�"�9mZ�W���<c"�j/���5�a�
s�>���+6�1�.�z=y�*R��
)M/?o5�G<�J_T,~�Q��b�>����a�;1kE��_Ŵ��G_k�o�xB�R:g�Hy� 
��C^��F8X�j�3�:���O[��F���c`Ia� v�ϓ��4+z�Ng���E}#�uOW��b���j�OO��"���r{y��c- �E$��9��۔ѵ)L�ѵA\ ���C���rA�A��r&�}r��O�5M�\m�������ު!e�xd��\�	<�hK)�"��ta�����ֽ2�^�@�!�rkR}���V֥	�t�8z}a1�K9[�n'�>?���FC>^wH?|ޭ�M̈́"��tq���B�E��.t�\�q����4���w���#�#} �����E��Q�y��rF�?{W�Ӷ�E9㏇<ۤ��˦`WXr�I rpB��(�@i��i(�U�������={s�x�yi�Uy���>k�%ڢ(!��eP`�Ӯ;��K0qX)�����9
tB�_x�jr�/S�tx���ݣ@/@Y&����l�C��'*YS��͸�zڌ>4�ab}}s���-��0b��.񹰝�l���*յgx�:ή(s:\���Ӥ�r#T�O���0н�h?l�'(ٜ-۹�+L�A֕j��O��P�St'����t:��uA��}M�}�����{���*��Cafg�h\t]��#�1�h2��!!x5Q~� $���k*\�Y�wH5�$��(a�c��Ү;we�f���_�}ۥNz���o9vOe'�r\\����.��N�]�Z�����u�+����}��6�+Fծ��R]8j���ݖa�o
bV�&�����o�F]fĆ������9@����]\� �������~��~]�3h��n?��Ư�I�\5�"JRI��9H���/	�2�����սl��j�p��k�n �G�D���QR�t��w�sL�ϯv:�j�h�ϩ�g�����B�9P�%
t��߀��C�@�A���˧T�,���?)����O��0����''�e]�Xb݀̂����V{��`WiW5����z�@_0ꦍ
tp��mUE��91g�T�Kr�M}@D�ʐN��̹�����^�6�~�Ɩm
����/7;+��EQ���C-L� �Sze�G�q�Rn�^���t�����q.ØjoHf}    IDAT�ђ	W�eJ����d֘]������m���E�u��:��$�H��Y�S�1������5�ݴ�W�"ꕌ�(�� f��!$�"�^D����S�g̫��)�	˟���"��9����KKz!o��k��/	�o�֓�ngL;3����Iׇ庡�)��&7�ݲ)M��tzS����h�SjM�,HC�Ai�F�K��988�� ����������Z;pS�����%��-P`=�؅�r�d|��Z�2�G6o&��ݾO�g�A��N�q���F�)Sݞ��Ń�F�8�]r0^4i������6v&��6O�n-޻�&�dEJ�TN*�ok�RR�G/���ܿ�����~j��6��,�nqq�[�s�Uh�QF_�b\��J� gLQ
���z�CY���J}i�������S�N���\�]�w�4ˢjWdQ��%hƭu~��bG�d�N���DJ�^Ls��9��ȉ�ǡ|Ouw�q�<�d�$E�Li���=ӾAq�M!"��������2����_G�NwS�,�l��)D�f �]��4ͳ4*�5��@������vg:�8wq�f�]��jpS��J.�T��\a�8D.�0<�����n�����?����s�
�
��w�:~{{��0C�=��3� )�j�ڇg7m����o���/릨s���ޛu�)�J��(K�hחs�훫�8r�/��ਪ��k����O釪�Q�k�P9cd޺ӍI#���1Ǖ�����*����(�m���@����f����ҋ�wݏ.����C@wVi8��u�3��S����\$��� �����c��J����|�<��V%�Ⱥ���������H�q`���/����?��j�1�v���J}`��R*���K�|����4\C3�}�`A�����|=i���u]�۲T>�N-��!Ϙ�j3fմ�s�vk4�\�Tx�L�������uU8�hN7�Uׂa)Dᦊ@x��B��*�^�4�9$%�����[���S�/�\;ε��3�8n�Љ�]��&������4CC#"���y>==���~ �(�T��jtdt��Რ��,U�"m��_{�{��L)M�+������.e�Mzq�T|�G��}�˺�,K����=c� ��!ga��HU����9�
wi�;_O�]Q����Y�L^o	��.��"��B^h���@d�(
�K'�(�1���i��rv�]
M}�̲�8(�ۍV�ey��?'冇)t���t^E嚭��Px� G��:�QD��N��6���I���uOMt_N乞x>s�����L�� � YHJ�t���g�+fҼ9���R�e1<.����?�sD:��"�vi���+E�.Bv�����:�pݏ��bLU�):<hǔ��ͅ�ޗ�鿼^>�?|����8P`%����6��,dDŖ$��j>G��=:U����E��4*g��qB���R�����w��`0�o��+P���V�	t@wL���j�D�cĞ�Z��3J㞣�w�h��}t����uz��8�4UF��=��!{�A�� >}��S��@�f��4*��A�I
m�V�����פI�}8�e�Z�K��k����(�a�1yzƆ�rn��t��+��5����T�=��/萙4
2v7J�χ�f
��>�<���)�q�`����f�2:��dQ�A�����f��j�+���piQ��WC�ݱbK��3����.��	g�3����޶m�C��8`p��u�s�S>�}7&�ϼ8v!I[S!�F!KEu0�hO(�W�� H�e��Cr�޸�\H��cr9	�L��WsYlhTq���yV����vX;�d$�����g��������SMj�����WV��%~��������l.˅��w�?m+Y\��~h�P�p+,Ңdk��I��;�5��DI!��j�QHi!l��^D��?{�o&iw�܏|�!���A��<f�9
��.��!�'$-�����zH}-��61��%�������"K����66̐螫�7H'_YG����u�tr�e`3}���"�6!"�iFW��_�,V��BG/xC���d����z#dr]����-D�Ɂ	gX�㚳(��*҉��q�	�V-dGo������Ñ �"�Z��нb�]b�ԙ�&��c,x��Jɩ���.��L΁��17�qz�:�ꌟc�,bC���Vw-�)p_#�Ce�Y�[�7�u;�����꾠�ݗcpHg:�q��躨�^	�+Wן���.�$�f�-����g�:�#�����$T���s9z �ZCភ�k�ޢ�-�%,���,�l��53��)f�<ʹg��,>!\\�g��d�7�W�B�u�x g��S��`Qx�F6�+����~���j��>n��4nH���'G'8�q���ϫ�ə�
��:���ǜ��֠�k1��DAQ��.��v3��"�[�G_�C}M�1����cy�࣋H����1�lO��v��4sȊL(��r��a�ДYA"U�v��*����"
��i(X�&���.�X�¾�FcIX���)��G�nQ�p����l�;�-�3}Rp{�^��È����a�ɱ�j4�^��K�, :Lau�,˪��q�"I�/�����������,[r�;���<#���uN_�h��.#h�y�zbi�""ߧ�*	=�,D�=�1n˖%)aЉ�7It��!�R�1�z�����H���	^�4iYLް)F3�u�Q���/�X��r#�z�'
�#x��-���]��X�C+��Ѳ!=KZ5|Nٜ`!���$^�m�3]dq��,
줗7�v�yg�`�L���`��t �[+|B�\ 
lyYS	��"h����Y�O潶��C8��0����/ol�qe}��om"b�c!�a�X����B�-}�zJ_[ }A	�%�(��8����W�Ÿ�b��I�^�Va�8��5!��Mx���LɔЃ�,�&�kz�������#=!���M�!G:&<Cu�&!C�fs�p��=��k�.O�ȜZX�g�z{����nA��Lo c��)L6aT٩�=�W%���ܫ�l�*+�,�_b�t�σ�ı!�'7�~l�;�/69�ۘ���m�R������ђ�R��b$j�,JO	襂���&��A[��z`���2��^~������y������(�F'Q1�O�xE��h5����0�X��d8eg��d����'��-2�üg�8��t5���ۥg�j���i`�bqX�?`�j1�7��<�5���ӈ������3��_n�H��qs���
�$�[֣l�UWe*_��Q>��&�����궄@�"��*�{\�<j���w��Δo0o��i����Y[�x�������}<�y��1.�h��5	�k�=a���Z���V�%M�uA">�O0�0�{�$����N)�U~��A�����>�3�qԽy���j������ݽ�7u.�ۆm;�>(x������o�����^��=kv�.ϩ����)"��roZ6^�
�Nݵ]*"�{���4}��#ˢV�;m@�o��Hl�N{W�a��?I��qsRՕ���������/f����wP�5��s�NɈ�J),^��x��k�S}9�)��E��?߂����@�^z���J�˲��il��8�[��v�u�������w�p(����8�m�nz�<�u�'U-/l��,�1����ǝ7�}N�����y4[�.�v[��.������m������xaعL��X̐EC�K�L,�Я����rҟ�\�]�q=�&t�߯y��?���n���"�������뛛�������#��=;��F1?�~��o�x}�vv������L#
�7T$�G��J��R$USeyὶ���ѷ4M2l���R)�JۗeC���bG���v�2��0,x�a��p�rq�����(�1u��=��~D��.��kvz��)�t��h�a�n�)�tȪ�| :�_�����}s�<e�(�S�Bz?H�����쥈Ԅb���$<��Z�ժ���'/qϤ�����x���}}���ER��9p;g7��Ӭ��4�ίN����LT���J���rKT�|��� *������o�����;i���6(����jB&�(�H����7K[[�nۊN���L�H������~t��b{���ZT�۳�YA���-�:4 ��(ժ��Þ~ ��|8>2�m��������u�yP�i,Q�c]:�m��O�K������o�<Ǫ�"�f�Λz̈�d%���r���Z����t4��>�F?Z��op�������}#M�9=�� ��W���R��+/�	E�}A�Mx�I�b���D�Wu��ɈK�`hL[����+���͠��'�F?�tX9�o������%Y�EY@���t���f��`g�$k�������6�#a���㠃DG�u�o��xP;0?d}Ȃ����0y�l�39�̰0�.����R{����J�[�V�v�W�U�T������7ш�%���'��aYKv��k(T��A��q4������j�v��\����������o+�R}�����>���.�h��w�bG�է�^^\\�~q����g�}��ӏ'lO�?}�B��O_�P��������>���8o�*+qR���X���7�!��P����֕��ǑC(eb��U}�2���������fs�����P6ܸ��n6�t�n�v��>v˥,�]f��������Ö��Ղ!��u}����{s����'���FT�y�e%��EjKZ��l�4�n�s�l>��N��(��c:�K�� }������W߯o��J�u[M��J2�׳�����?OnON��n�v���/�./����������_/o�u{�rv{r��ER�0�|�����n�o9��Ι�θ��F��E,9�<{|�^�9�g��Rv�aEf���B0�~u���W��|�3���c0��s�T~�X.�>t��w���s��;�rgk�g2u���u:(���[��\�+�7��_�T讒�V�����dO�H��}��[�J��^r�+���-�����n�ۭ���:Ξ�9wG>Ga9�+��[��������L2���θT4Q���OOΎ��,9�e]��{���Xλ]��nG�d�wt�宓T%�P;�����]JF)��9Z�D�4I�)�:ttg��
C���tYR+6Bg�$0�aTi�BtZo�#1d��&~�^�Čf�M�6���T�%zr�y��-|q����/'�z<MF��|<�F��d>��g#j͎�c�>�j��rFW'���h4ZΛLO۶��!,h���������ӫ�פ����qC9,u_�d�O.�~��!��ǔX���ʍ%��xIp$�q��6��U��t� 8G���t8h�h�6���o����c-,�cf�*
M����*���q�A�5+�s�y�b��9���3�LtCp:%YB\d�J�y�����G��O�yË��5td��XG��S-" ~@}� /JTeM���AēA�͘��X��n�����]�?9���,8O:=�����^w��S����)2�<,�lL҅�p�3f��Ɓb*�%���ä��73M��$�����8�y�j���������y�����������)텶�ǔU��g��o��'��WHdi��x�Ś�1GP'D�[)Iv���d�Ӓt:;G�m`�c1�"���5A����L��ȻL�`��!��"�����	)�	C����F�E���'x�;���IV&�KUW�P��\�W���=�Y|��֬xA���-�	X�i�j}�^�`��\G?¤Z���L�\;0pb�M�Ip�ݺ*&�-�DP��0�mt�6Zj�b�O�T�b�aC�W!�SK@@1����9�;�E��Ǌ�zHB<A�˦�Bgel&.���^͌I���C(��X��T
A��H���?.���%{yKl�6:#Wy�$)�ʥ�bW�X�h�OhW}f4�����G,GzyQ9B���G�������������R�h́,~d{u���6�Դ�N����amvpEh�o$@�k|�{ 8�E�h�1H7g�P�~4à�����9�c��S ���Í
�G"&��0��n�|x�e���%�/��P��gd�f�킨;�C"��[^1b5?lc��fe���*r��������r�Y��Y�5���L���mt^%'�,��9������3�ɳx?L�7��$ �$ �v�\�5�0]YoY
!�!�N�<"����d*J����CXR��DPx�Z/ �  �c��o��� x�.�3�Q1�Ad@��C�#�*��xG�R�I��-i�?�T#��(?��R��Jqi�^wP�B�p��m���
X��*�(r���gV7���������'���v��,`�Wv^����Y՜�)ُ�7�a�c-�t�|�Z�x��X|�	�P��s/,l#1@R�h��zO2b
�<�x�$4B�HRÎb�(Ά�1��Z�< l����W��5�DW X��u��~;�:=>~u5ׁ(�Kf�������>-)Ƅl�x�~�@'�����]Us�9ø!5������UUղ����q�R��y���S@��R96
z�������l�g��į�@���R�ȴ�0�uv���{�� �ĳ$8��������kfE�(�3 t�>���	P�NX2����uR�A1sW!V���!�`��钵 ������X2�ag�O���Oh�i��@ǒ�/����{�p��)�^�n��oB�*XS.׋ʜS�Fy)�yNWר����^d'];q�R�Ħ��5�tЂ�/,?��':O���w��*44��_���$�3-��jó�eI,U2�Qx�5%E�(R��$B�0GT�����P��Mq�=�f:l��8���ζj��hj�
��!5�筭"Q����@�;�{3��j�&z�6��b �Pt��ŤR�8��㲨D��_
��cꔼ�L������O��dB�f:�6͔'�t�I7�,��|:����x6M�"���w�Q	x:;�{�ڛ8�E��ؠ�W
Y�d�	�!HC �'&��a+�		d�,Q�l�"Q�!2��d╘��{O���]i�c>Q~�u�\6��ު�XZ���IS�L"I�"R(#ţ�P������d�I|!��;H]V ���!�: ��!��#�/��W��"�U��oPUܲJ=��j�~$aXF�B»�
u��%J�Lr73��ֆ�s��::vC1d$��D#����EY&	�=	�	`����@=�Zr����Z�@_�zڈ@D0
�J�Zl�J$�cE(X�$L~qV�  ���	$w)XP�&R��&^70L��ɾ��������"�%6�<�f�7���K�'L&a��e&�tZ"�O��)
%�-��J�WI�-�^+���=�NH�0������b�+�Q+�Z�ε
�
%�j(��\I�zH���x4��;�,�2��ξ�����,|-�J
��-�D�|TB�Q�X��䐀�5��=!���/�˲�4��dA�k�AF�E�|��RH�ڨg9�U̙�CL��"l�wM�'ڴ�U���ص,w��ϙ�����ʧ�0{Q�Xb����ɮi�v{���]sJD�7=<��@ �����[�c�r9I�bL"�z��\P��qy~q~	C�����\r��"A�*���0c4�c��l��ca��
cW'���?��}�}�?��>:�L�=��F��+���U�1CW�q��w)*�b�X(�k�$�'��
�ؿ �"�(�k�A.���{z�|_���Fx&��*OL�����-��j��k��kۭr�n�� @@���6Zp�p�ݖ�p��p��;Ì� I<&b�-I8�h6�&��Ѣqح&��8�2�)��l��uӾ(1����"�$s��t��V���D��f��)?�MWy��j�ׁ9+����>#�\�HP	)"V�E]gW����S��������`{��P��>l��V��������ꫫ�Ց�ۮ׏V��?^�,�iy֣\�G��C!��Y�%b�$Y��a��[�K'iC�$e�=�ֈ�5� �!�BDPY�͢4J��    IDATU�0����X�ܳ/����GûU�,�$���<T�I��x���?�������9��sk^b�Vpx�=���"�wDxi"I�M�A��U}���o�L��Z��ҷx#h��8�4�1]�7Ln�M��a��<u����3��v(�t����b��(���o�F�q	1�D	�(�U��w�`�Ӣ�̡��/��H/�uY�#����r�x�zW�E�F�d�4.�3��`jiDw���,��s�L��,���'�q|*v�q�=ǧ�p��pLs`�&z�ދ �;�@��v]�v���E��|��>��^��o7 ����.�Ωe��$��5K��.��hR͔�A.繧�#H�<P�!Y�|�z? y�Ѝ6-�HB��n���v���p<Q�0T�2;�p:v*�����5�k@����8�#@!/��A�������ScК�F�LzZ��zKQ@���d�"��!�:�])��QM1�{s�
�*;�p���]�+��7��_���{���>�j��/�,Ft�Է]�s�Ο}����[:����-σ3ݠ#���mB�����:� JI�]��6���GF4e|�o��6H���c�+����L_�Q�����Q�#O>v@�����:���yx���Ð.O?�h�s'����<����G�Iφ�{&�%����'�EzA�/�jL'�{�y�tY�PP�W�i˞��Y�n���k���l�>��3v������n��3����f�v�n<{���_j�sN�T,ʓ�nZ��񌞝͸�3����9���p?���Y{w�tc��m?W��C��a�(}k��rsU�������7g��,�ngi�>K����Ym3���K�S�7�cV�WL%��-J8�DX������?O���D?���������z��f�����!�W�l�t����u��]q]]���{��UY����}��^�t�$�hL	�C&Y�����X�ɧ�k���EC��T�dA��T*�����m�WL�KN�&�ŦA4U���n���IK-穑eM��k�)�Z�+!�J�F�W�i���m�t�~I�b�c����{;g9���m!^˦�i��V���mmnnm�{Q��@O�7�zɠ�*rkQ\R���ӏ������_���(F������S!!�'�G��Dh�@3�X��	��.�X̺/ҋ�d�rLL�j���U�]IE��#�_Cb����f��Y>��i<�!x-���A|&�v-��Z^Ni)DlBW�h�����Ӯ��^Sú@cz,�
�ɴbuog�D\B`��얶k)mym��;Yf�#����P���7�7�e6G5U�V��Эb��!�*�/�At8������GTEzc���j�l��6v��RTx��M����?�~~���덍W+��++����<�a���o�W��o�ol �⫕������_�]kO�ZU&������s�ˆ�ŚĀC i䐄��zAe(���.Q	"z�[��?{�:��>�4@��'n�:k��}�:>�-[��URN��Y�`d�wVkK����3��£���ҽŪ.)�/��׆g��x�Ȳ)j"����t�7�ݿ�^=�Y�S9!l|��
�b�tWu�A�0�'?���{��%cIV���^w�&ԅ��@r��;��R�:@�`t|�W��_=��6���&IlG�#ᷰ�]{��r�)zt}'�2�':xj�vd�컀��
�6�oz;���!��:{F�i��u<��K�j�"L���J�N�;_vr�R��+�:�jυ1����Z}�c��x�pNf$���@{�Hf�
_#�krZ�΀>���]�f����x�l��6ʉ���%�����`�SE��+4'�Up�=_�|����kю�����'O+����k�mRX���n�vu3�#�E*i���,�g����-3[�����wwr�{n�?XϪ�(�i��};c���+ ���"��p A<>�׽�'�O7��`.A-�~�`���� =rLn��\��>�W#s�R�y���W�ȯ~���Ǉ���\���x�"��������BF���P�����^ ��wOj5>�����z�]��ٸn��GB��
ȗ��]P�Oh���I	 m~H8��	�{{�s.�+���e���A�M���!U�h�B]`b.�[pQ@rw��`����;�p��%Y2�HɱTJZ�4$�'�/`�?������h����z	n,K~��!l }:,,fS1����]h����>ϕ����\��%������2ׂ���c�����=Ϧ5RZ�X#q��R��e�O�3���+2:���24�o�����z�5�R�%&i4g��`t0e`��
��g��m��!3^9�ʕ��|��6��O�A{�����T�� ��N>�Y@����b��uEl]qL�U�뺭pj����1�w����F2%�F@ hM����]F�uF�#<K	t�� �_wm�u1I�S<���!x�>�C����D�.��G:A�@rI�%��q �R��2����k�m�/�Z^Nɋ����W9_��oo��q�Lkn����@ײ	C�
,�3 ~��n�g��i���%�,�
�9�[ۮ�}m��D@��������;�����|�������&��B��k_�b��i\�[���V]U�ܙ���b��v*S%r=���K�:�c�vP	#%�S�O����x�����X���X4,�p�#M�O��A����ve���D��j��ã��m��!ߡۡ��U�FN���/N'�s�^�6	���B��q�z:͞����KK;�Ť��[r~>;����Wz�� =�5Зֆw�MD�l���F\���۞n߇n����r�UUpt��o�.��$�f�	c����t��sk����<��\׆���eG92ǴM����kt�֔�ϕC�t����e�y��O���	�6r���������H�E��^WqU�����e��QW�W�Yfݧ���"v"���[�btBWx�W����Q�����W"NϕI�D:�����	b��`!Ǥ��>���龘OIE���}6^��sC�6��Қ��VL�т��]��]�پ�1 ':���I�T�O�9���C��u�4M0���1��ӷ��\�4#����x���Q�k��;h�g��/�׵ ��X9�骪�޷M1��Eҝ�� �Y��F�Ox;@�|�E��x���'�3���Bܫ�r�o��q���%�`u 1������J�r+W:����)���v��}�R��;�uB��/N	tv�bYm2ɢ��fݗA�R*�����g���熖5�qI��l�l�U��X�n*�d��5��v���έ�U��n��m���#��L���KWwMӮ�-�6�;��7�ؓ-���t{�^�y�t��3���T��'�?��g2��R9��g��C��q�@?��"G9����j7c0:�z�rG7ٰ<8:��C<�ṉ٨9 st,
/7��^{9�J��D^.&D��ҽ#2qe��R��٬������t�}��+�Ky�e�J�~���C2z1��bVnb�f
�����̼��A��|��o�l���"�=Jܦ�V��C��$#���.E特ý������iz]�mEeX��U�'�n76�ܜ[�g+���v��]0:�{��'J�����N�ݽE��W/Cl[�n7��U���=n�B�Ǚ�bꈹG������.%�D,�J�S����1:>���Q�P7Gw�s��0P��?w\\o��{����]H�"[G��<�qG'G�}WW�eh�\�r��?���ۗ�/�|��_o��q�	_�V�B�瘔/��/� t���Dz��L��N���|+��f�Mv��x�ݐdYk��[T0��$�m��R��8�	�[.+bBGd����dt����l�}�rs��9+��X��w��yh�L���Ӄ~{��kx��1�g����^����puu����t?^���{������C��rOH���.֦�ٞ���)��Rk��b�ën.'p���=��y..۟}?ϋ�_�'� s�v���}����l*��-�Aȏ�<�>��gs�y>��W?46w'�c½hZE�ER� /޹}|t�0�B�q�,"�@����N�i0ng��-/cc�^�U��g��B鈽����_��_�C_��h�mV=��t;�ŽF0��s�ѹL&����D�M��G�xL����/��}���}��Tic���\�l���2�xey�;F-����8R� ��^�:�_B?�ˣHql�4��"t�����n-���|��I�3�^��2��@��t������w'~A��8-_75�.���v�W��3����f3Ө;�?�c���QA�;�Gϟ��2}��S�;�XGW�G���R	��2�������_?�@����oc@�h|4����������j.7?%�g����|�,I6�"�M���:��3R��1�>�� ��mH�Z�'�k�n��M5�Mɍ`�R�4�7Q0c|�[C�+�x],+����㠃���B����;��.�1�=����*]��cE1� Qn��bAwH��c�<��<"�0l�����65�1I(�ͮ��{u:m��;�5,�G��ɣH�A�� :�`�p4���/��h��x��S�QX,����A�j	85��9u������14q󨐩��9�?==}����?	�G���(�G����ɣ��|!+�h��3�u4�V?�۹[^!����lv���dt }C�U�љt��n�l� �)qy��v����m�u�h&a�Ys�Qu����M�� ��gAqT�Z}8����鮗X��3qb��I܏$|���"lQ���;��]���Y�ٳl�d}G����q��4���F��yu�?n�<z��@�����$��ncg�5FQ'�F��o5��U��`�S�Ys�����$�d��������I�[��ԧŮ��G�����ܼ�m���0~�wP_]̡�|㾜l.ɘ<�%x��!������2I̝�����@�#E�sys��T+r�'���&��ڍ�'��Dn�$�u���'&9k��`�<z���6m�0��QOn5�ѷ�WKy��y9��髡��� �	��M��[��^�7H�G�MoSQ4MED�X[ם�16-��?�ۅ��;�J�X$��ݼv������ʓ�{ݡGң�p�舺��by,�Ya�ߵ�h������8�}����^{��'�~�}.$ߧ����__��0�mc��[������.�y)�Y�U���˝�t@�"�����ϵ������Dq����y��{������j�I��Rl��m�=0�(B7��,	�!u��c�E�Nҝ�6%�Ua)]�٭]�Q�f�vG��R!Fw�)�Ѵ����J����X��O�f�� =�܌Ζ>T?�������"�f%�1���^��/�;h�'v/�}ϷM\1��:eJ�1<:�y�u"&��*�,�
&g4=���yA@8;�O����a� �����i��m}^��,����$ֹH|�S�M�I�+�T6�_Z�1��h0N�d���tn��X2��\:�E�\~����
zFuG@I� ���O�V��H �z�X^7N�(�������q,P�f4�Kj߫�ȣ��"�  tyXѭ����rC(̒��<IwD񛽝	J`1ڝ�d�Yeyt0:���v-o�+:�e?t�D�����F���+��;vs��w�c	N���!Ks��ޝ�{z��E��ș�� �uyv���s��ipn�+�E�`��ߏN�xE@��|�^ȯ��rf}�M�u�^�d�=��}v^����O�$���ۭ�ՍJ� $s��4_;'���5-��K�)(���Ehct?����b٬��!1�������WWyl)'1D:�M��`\I�!�G ��޹u}/��:Iv32u]Gǌ^4H�k��d�xt̞W��$��2R�Տ��n�{��EM11ZF��j�\��	1����b��_�SG<e��@���};%�L;S�*��/��{�,��zX��K�]�)'��rS�>�zF_�������,��pB��!e���K��R������YȬ����$�>c��yY�.��%)�},XSKK��4�tX\%��M�^C�
�V���E��O����~g0�򨣓��Y���J��w��+�T̥���B0nwi�\�5��4ù�]��gw�ޭ����R���ME0t�0,��=���5>������ֽ����v^t�Њ���w�#�/�ߡ��(�K�Sb@���IlZ��k��g�v5��*���9���3�y�X}���I��
����o��<:[���Y�
I��Va%�q��,I+3�����C)K�1/-|�{�M;�9��-��QE�~��a@�"����l�b�$�bE��Nv�Vg���щ8Y.�Fg��_��x&��r2�:.������I|/��hCe�BQ��h����w��i�YTd�������X8v7V	/����8f2��V�M�M;uK@�Z��&!--�ҟ��<d���ē(R^�����{�=�\Ϝ�C#�������O>�U։�wP��j�l6ΥGo�v�
���Aۢ'[xyS�;x?	��t썧+��`c�UD~�aU���eU�����(�7	�/_��2��}���<3��8����+�������j���L�>�_ :v�?O'�$v=m�v*����X�(IM)�T�-�]rtY��</S�^�T~�÷���w"�n�i�.]�A��I���2��I��ĮG�i)F�{I\�/�Fg؊��KC�b��z�8ze�%�Q`-@�.����p4�׆#|�mg2�G�K�1Ղ��3"�.���Ou�q�8z����˦�ʊ��Aی���`�� ��C�~bC�{b+'��A�R���c�#���D�_��o܊`؋�y��?��?===�/_.�Ο@�^,7�l��q��/��{-�˥Q�.Ye��>>H��ѓ�dv	��;���jSjb�x�Rw���y�� �ʸ�w.�aV�BeL��9�uʵ'H�G��X�S脾T�:]Q�9���Zg���
�'`���J���@
�h�5Ot�":=p�Z-����?MB����B��U��:Ο�l�#��1z���[{��GEц3]6�T4c\�+c0n{ts=�;���'��n�(���{�k���q5�.����C �ͤ�Ij�o����|�___�{�/��a1�4�n9:�qX��Ylq\y]۬<��N�s<%>�����%G�K��$�\y���v3&�%�جB����y���VƠ�B{�
ttּZYf4�AuF��(*��n1��f4c##D���%At�����xԅ����2&�4#��<��N'g�������L��j�]�i�w��W�j��S�8A���%����`ڼV`ZF��/p��;�f.=����Q��63��-{�w�<���ݐH$�k�P꾐�n�Z�,�o��S�^?�@��t��Ki��F�Xd���Ͻ�P�Iب��Z�n��f>&���q����s�U��\�K�ds�y�Q�^�M��f��Et�� �7�`3D+���q����1�pT����4+��2s�$�O�t|_�R��D�@o�5�'�OC��꙲FIB��DJ������(
��8D�	aؤ�1s�yWE������w�n�3�o�隨&����p'�;�����YdRҎ�<aM6�מm�R\�&x!+�k��}���b>��<�v��Ź����uux���a=����,eʱ�N�<��s1�CVf�ރ$�.P"�K�/���[��������~la�j��%$S�~�.��x���Qb^��>m{~o5
�b��S��"�R[g*6��ڥ??�ʄr	B}��"�pt,*%��A�mE)e0���i;V��Z8i�^@�T���f����x"���dRH!���<��Ύ�Qn�O����	��:fYVx�����Ƅ������^�a��rBL�����Y꾺P͠G@���{��w���0���Z�J����/���<���`�U_;��ki���$g�?-�~�s�@o�9�sR�z�V+�^�]"�r28:�����8]��	�u����:qt FR�]0@=S6���e�s���XڨbR�Z��7���ĥm]"Eu�wm    IDATE��&����ކ帞?�kzS2�~XtP�vѽ��R.���a8Y���� �v15<L�7/���-�|�8�z�x4ǥb���r��W��_ |a<A��������Wה�?�}Z=��ȳ���7�p�Y{-�g����'�m?�����Z��P.'e��X����.Sw)!˼$o�{V���{G�'TBd
	�Z�)��BY�"��V��mx,���"z�F�t)�K8:dtb���C_]��kRH��$�^oG5���Q�D-��h&��c�3�b�]3��ۚU���mD�Wʟ�\;N���RNN�^�Q,��} �>%쑆�OD������$����ޝ7.��y�$x�		^Z�$�����؍�j�U���kVu�P��O����?�����1����W?�Y��$�e$�����676阌o)��|�-�]Ft��K<��Q�k�XW��86��v�ʢ��gC,ü�g�p4��ڄ�b�s��>�2�`�F�TD��*JwԸ���z��3S���q7[�.�8YP��$�ȵH0�XL�39Pۅ��1J�yB��m�LfL��aiG$#����g�X���9
�J�b��St`��ϛMB��~�-g2nvP��"�M-vB�[�/�!�9*.�$`����{���S��	�G��������j��C��e����ϱ���g�B���Z���L�y5A������<w��R\�g�[���?(u�I>��Ը�B{�Uݣ�f�d(�*��V�`B�w�����Z���O��"�2l>��{w����z<F�������r��X)�Es,��m��N����;Y;�@i�;Λ�tN�qO��^�ǘv�|l�@<=#�FD�;�0`0E| �\�s��f�)= .�5�%z��ίU�xJ.M�����������5���n7P��������k�iQ���!�1���XN(v���'�I�\H�fUZQ���K�P "�"ԅ$Z�t���3߸���b�
U-���盙���^���=;�}c��&��[2��Ox�N�]���@���޺'�$I�e�W֟/>~��QgtE 쮦��A�)�VBU)!Y*����>�9��i6iB��h�)�K�v�jL���ᤇS\�M2���ad�0q��$w��*��o���)� �<�����{���p\����FvGsG�5߄��::�'��[
S`���.{���l;������Q�QԞ�{
�qa!�I-0�cG�0��*�Z��}y���y�~{���q(��z�ߘ�~�Z�7�ט����m��]�e%cIF���T��YE�Q^���cvtO��нX�6�ʒe	($XHp��b��փ��'���W7=��X�h�Kl�vAc�L��{���JDI&8�	.��h���58���c�m��Fwэ���l@}���q��G<����!H�,��B�
�c�ʝ8�s'|�Џ P@�6���\����{Q̅�S���u�$�j����ۻU����ޏ�8�Ǆ�[�R���g��(��):�q��3u����-utj���<2XB*�ˏ-��뒡r ���Jj�<b��������򾴵�?��eAt��cC�<m�u�9Hp0����Z���;�
����6�i�6�4N�<�G{W�HC� �'=���k{���N�+lۣ�`�
!��p�Ҡn:�ɕ°2�ġ�4|S�{�ຣ�E�J
Ɍ����^�G$�o�;Z:p��r�@ғ�	+����N�o`��7��g�"^P6#�ڭ�~��u�)��Gt@w6�|�2�U���|��OQ�u�Į�^Rغ�{�ie�Ftj�"�
�q���_Һ^�U]ٕSQ��y܎��:�Sغ�G?R��$�wW,�ײ+��"s�q��		���v|���.�+��욾��O��C #X �hO�K��@���J>�Ņ~b���	��7���a� ���oVFa6Ӆ �	�I�����鎕� �%I���p�@<#|&�@k�9;�M<�<`���W�pGԂ[l��W� ���G�d�P���-~�E-��[f_�����P��ܾ�L3zw:��oty�/���6}��f�24��%)��.����O�����t_<�9�CI%#���}�^���(C�AEd�wNU��=��@#���Mvz����Eg�!}��c��e�c��q^�]]I�� �UI�Vm �'��� �(Pa�s.ve�=;\xԍ/[�0*Q���hJO;�ӻ��谀M$%�	ٗ��y����7ؽk��-����!�-�������� (�k���_W	]޾dP�[��?�^{���T�(��[���tA������f���z��/�O�h�4��֔2�ˏ|G�u�RԬ����x���Y3�G����|9+I,��0[+��w��!rU�:5X�6m�9��Fϸ3�>�0�O� /� �#`>\��Y
����U�jѬ�-4`�i,X�ݏ��`2a)���o2�0oEG��'�	X�'�����؜�t�L�I\MssÛ�(�zLꡟ8½���t;����q�A-��	���Q��u@�w�oݸ���ז���$n~���� ���ΟL�o����_]��굵��RGz��ygdQƹAf+�����Q��|{1�/�G,��]Y�e ֏ϩ�W���=�"�HjQ���G��H7r��6�M�Ӛ�4����B�t��Lr&+E�������טх+��X�o��>�;����s�Mu����A�_�`ѻn�Qآ��6�x0xs���b�	fV��-C��^N4�=s�R�л�!b��y8�����_n�4hL��s���f�j]UddΕC��}�W����+)�џ���D&P�n���u�ga��=ϋ_�g0�]Qt�G	UZ���X^�f]Od�ԋ��o�<^�o�5��ʻ�`%5���K�e�J]��d9u�ܻ\����:N�&D�HU5q�ꍩ��S�}?����ɬ���%���EEe�����6:�iB����Q�����,���u=!Po��������q"�Ԁ���>\�@'Sy�A�b:Y�Q�@0�����VxL��^�Y�Hjُ��83d��F&C��b������kkkq�C�G??��_<�Ϗ^A�r4sP߄ll�������غg2	�]��$�ø�BW�lҷ���/�ǅ�Y��U˸jd]Q�˒�� �����'�Z�>B�q�r�8��ph���wFaev�i��h���祝q�.��^~:�Y����Ĵ��lY�����D����|"+�v�s��w|Y�ݕ8�A\�m+g#���r4�� ����8ÛV��R�;a8B����	)�������^mcCUE���������YjL`�˸��i�\�)_��u4�v�N_��ȴ���:��է�LƠ��*ݠB��w�~QJ�EE�լ����-�G+�O��]Iҳ���O�VOH�L��PgЩf�O���z�	]�c�A�>C�@+P5{���Q��;�h�a�M�K`;�u�6
d(V2i�w�#��^"ti�I��0'x]!|�¨D�������w�?mcYT�-?�C>�	f�+I�#a�y@~5-k ))u����0��V!J3e�v;�KaV�?{�h��'?p�*��s�����5_&@�A3�2t���A�}o�s9$��`�B��d� ɨrP;���4�*6w��i ���z��-=G��9�	�f)���6Ly�t��8G�����o��}���/_����_�ma�KvI�U��9[o�Rl���E:4��~Ҋ��r�~��5?����-GdOo�mm��PES<O��>N�x'.��eY�+�Q!�0=ڿ�=:ڽ8��R����/C��|]��:�L!�9]Q3��N���� �˔����B�����Vs������!�M�g�g�3�'��v�w��w
�z�MÙ'D�P��X���y�$���ڿ>�h�(#2��&�_u+9a
C�s8�X��]�������g|eu��_��?�n���e�>C�����rqvQM�p���m��8�m�\
�t��-ݴ�%8G?8�*����޳�.�����]�z}g8D���^J�� !lK�e7_��gF������y�;~��EF�2
~S�t���{�~��C��|&��+�%_ѳB���!�|�n���3��(�b�/�������e���Q��|?*��>�����N�q�>o.!�Z\7�O1v���AΑ�i������{-9_H������������ju��soGt4�`�Ϲ�i�l��f2���9������O?~�'uw��r`�}��U� �6rJb��n���pr��8�#7b��R)���n�>��j2����1T��03y�:�ƞcB�J!��mtF�Y�	m�5��`����˓����ɤVdv0��Ĵ1 ۿhv��]!T*�Ɏn��?:L%�8Ç�$q}t��)��Pǟ�]���QX���ޏ��QD����U�����חOf��Je1�%֓!�/��5B�IV�1��ǏO�5��0�g��1X�*�I{�eZ��������!������3W�%����
u�D���5�W(D�8��9�JvQ�y)W�a�@�B?��]�rt5���Y��T��n&�e��
Q^�!���%̗��"/�1:�bM]�<:��]�h&�G��e6�u�A?�{J��3�i]�}-�������|����X֧�[�?�u�R���������\uO����"�a!DQ]]B�����Yn���#:Qw��ٖQ4M���%�A�QQ,[1l�,>O?~��)�7������6��ޘh{Ѵ��gL��r�<N�(QK	5g��(e���R'���@rci��Kd�_��}ݍ5:M
�����9z�z�F!���2���0�,����ŰZ�@>�%֪��$�^�t^�6Yu�I����KlCl�@߁�u���S�t��*���2�,��&��OcJXt�`�S�u֠0�r�Ű_�gK�]z�rK3_�*�v$�����rt�v�pnc"�r�dL�¹aZ�?��tͳ�4t
���)��ͦ��0$���ak�3�@�]�yb\�N,������%%m�%�t(G�th?	��:<ꌮ��y)0A�Lܕq��6|�˙�K�6��w)���E�"�٦�F-*�!��"T`�pr�����CD��#�/��(��>��؄|�`L������\�b�@{z��h�I�;�=3-����*w��1;��d9�y��?��k�VT�`c�s��Zqr����=]�:Qw�k��"��Q��X�rJDݷщj����XR��Gh;�Oz�(�(�G�L�����J�M�o�ϣ����T󈸗��r��Ǒ���|�F�K�s0y��9���-�$�-q��]V��$>&6@܂�݉X�ep�.�
@�L|ه{�K���������8�)���+֊=`z-	�I�mu!�xO�b9���=�U������M��Q�(P�� �_<�juϬ�Ė�e�RꞮ��LU�t"���|Zkb�6���RU�?�v^�8^"Ds�E����NX�ɉB=�r�����~��h_���'2�w����}��y�CL��N�?H5A�x;]!J��t��r��+�8B�<4o*��n��� ����[�
���J
�u���6�-M��~�2YGS��[�+��18ܟ�?<,'�l���ob~�n���0Y,���*�.��am����ݶ��TJ*]�[��:���c[X��j�hv��9�st&�\�"E� N~��=�~ɟ�z����;��+�P-�kh�ר4�������_��10M�9�/����rQ��<���{w��q�n��Y$���Z�3�u�x��X�P�EϠ+Fl��Jqn_�����Eð(kYo0�x������Y�p?�ʢ�� :2�j��d��<wƽ9>K��rD9T]���b�0�6*6j�����/]���x�3;Gy������3g��|���Z�pgȈ�>�A�����B=��(��hu�^6���#S�&$[�ˢ�}p=EV�í>�d|m���Q(GH&�8�N/v��h1�Z����A֒*m9L>�+�� Xcސ���n������T*��krQh�J��� ���W�ogS������_��oD��F���Eô�J��Ow�3.�X²̢�M#z������e	��3YV/�V�ƼmUh�e��~�֒�,[��
]��{+����7W"R>`m�oH&%|���@�B`ӤI�7AiNWJ�����7�����}���9眱�ό�3C�EQ�g��b�j�<�����$:_��W���?�dSht������s��Y��J���C��$������c-�����kX���\{���:��_�M���CO�q'���l�P���'ᥭ�Z��j!��
�sFjF$˻%
�h/ZD�d�-�Z��#���u��y���Q�H\���9��~m���`���IN�#n '��A��O�b7����`�<�DWtAV�{�]�`�ʲ.pi����X	���I�<)�"�w'�����a���|5������c��LiR��6/-����"ۣ*��p�骛��/��zy��f�O�?�S���&�&We�txU^�=,�^a�y�}ݰu҇�2}�����z�q��.�_��VqYe"��N5��!I��u��������	����SM�i���i�]�F��cco�����yooo	�����1�K�?3��KǄ8�;f�{�6�����3YHp�%#��v��JUr|���ҕ��'�xN��'tӌ(��5������E$H��T�E)��
��T�w�,7��Ԥ���Q���a>_���9�Wr�ә�
Ǿ���/J�z@��2��T\�����b���c�t4��.�L`ӗ��
r����������s6s����w�e�fŅ���sb���q��%�S����]�����׿~}l@r�h<�P��^�A	�A���B���m�6�5-!��@����$����iSa�g���S�<#�/g�ԥ��Tw��I��$z��i$�$S=�ԪN���`Y/����)m[��P,f\׵��2ۖ���r����y�ʥ�6Uf?=�����N?uFU������p�
��X�
�Z���ӵ[st�͸��w{͝�:�a��=줼 �+��J�ݮ�*8hAŭ�j����j�����R��uۗ��*NP�7;��k� p�\��]ݵ;V������Nk�����S����=�Z��GB��-�S��^�
��G��eȿ�t����	�1�SD1.JJ6�x�����٬����HW��=u�9M��&j2={���ۧj@��� 9A��y��,�
6����Q�����<�Q�4��yS5�l	
Z��r�a��#p��*ǡ�\�n{�`p�E��n
</���6�5��|.����'�� ]��=�R���A��N��f�0U�'ӷ���9(�j��ݝ�����m���v�v��j��Q�N[V�m�ƨ�,W�-��zv�ϭ�%!07�+2���vK[[픙�$�:D�ʂ���N�E]�k���ˢ6'�̜hP�E3i:��W�z����!��AФD���m��M�'o����rԐ��m<u29�Md���t�Z�!��e:=�7��`�eC"O�.��b*�McW�m�z�A�^� ����s�9������"�`�$�:������5�?�s���a�{׿����N[S��g����[@�b�������s�&h�;[���l�ޏA�tÔbUk+��x�IA������B��)t�� �0P�i�:l��Խ�m���T��N��S�V�����	r_��3��yBd��R��:�^��v��7l���e>����
3�X/��%����z�T�n��Y��� I@��N�5M�&Tb<=C��dEP�j�t��=���g�v�?��~�~��*�����)�� D��u�V�m��>$�;��$�0��c:�^��8G������o`���+��^�-KJ�'��2/D�5�6N�'�~w8"w�����?<9��7T��Lm�S��@Q!d��$�n�a��gk��v�H8�0 �`̓nؼIC�GyÐ��.�`���    IDAT)�:���m������^���������9MF����M����~��"�2cRA�o��S�]W�P�U騎�F��Qu4��Fg�(5J����,�<U�RG�wj��4�P�!�E�K�o.��%o��C�pCIdW�������n9+:��do����!%8���Itx#j��̨o�?5!�A�x��9�E��S7M?����j�Q��Y��9�E]�ɟ�(��+��(�J���lꏄ��ꇡ���Ԩ!Ȳ��*%9�g�	.��
����d,�Nǒ�$���r����4z�@��/�1Up�P�゜�!G�vŦ@8�ܻ�$ʲ�H����ﷀ�豬Λ�3yM��S>�h��<�H@+�x#�H�B�7�Ftj̀�27pSc�O�a� :5	=bʈ��(O�ǥ�:��X�a�q�S�h�c6��'�K�ف�)��J%rG���L~Qo"]��%��֡c�75(��c��yɕ �h b�1�2%������=�KV���Ȇ�2����½������EC��h>8���n6�W��m��*O��3gA��P��NY	�)�����ʦ[��f�u[e�Jm�~���v����)��>m���{�P���ˡ�Y�9���ЗvGFgX��F���.�i��5wY��T�:�j�u�2� ��u�><�R�-F`K�G�K�DA8GF�Ȃ��=���+���z#{��Jl��#���ȃ�������;��0��3^�j�6�'����0��wi��x�����π�md��T�8e|��F��3�U��s�&�Ķ6��V?0r${�
�����&>�×�B	̂ퟗ��������*�d����@���b��I$��A�o ' 	!SC.�QS�� 	�Az���*��%2��q�K� �s��|B��y��1ju�U X_ѻ����cϚW4B��X��xW49J숡��V���h���P��;X%�ߞ�a��Lρ����٥P,h^�Ś�x��N�\ʹG�8ۉfM�n�=@��]\vizZ�~K�c0�xɐ�͙����59Y�Xj���L\�0w���~�am8�W[��"MD�[k,i�v,gg��5�\�&��Im�e��O#���p< x%h;r���bm��v�p�Ma\Yh�ܬ�������jh��Vb�b�v�����;)"�'��;�4EΖʏ�͠�!�g���a w~��2*��G�r���R2��-�}i�dt�!%��.N�(�V���g���� ������F��P5C���<�w��QZ�Ȟ��`p��3�3@ETQ�eЕ�(���B�:T�u[K�x2��п�.
qכ���Q�+�r|�T8����șbcd�γ��wT���S�iPz�kgD��a\��ˮ_�� p'�ϬyX3�dg�ep��u_�l��Ӱ��/�~>�O�认\ ����>� ݙ k�̄v�萳�$�x蕄83%<j������U60jI�Q5��$�t8(�!�Qj�{"Z�5sءvm��(���kZ	���az�L,�pK�ӢpQ�
�4���;�T̰4;[�?߭��5ޗ��T��ɜ��zR�#������E9ޤ{n������w�$�0:I�Eݽ��t�]�CaV{Wʴ_���;JwHɩ@J���T�)�� ��8���V z�f�W7\)b��9�֋�.�R�3W���R�����e�����U��q�X��%oň��d|��ct�n㳸���U�]�U����.���;�-�e�@ˢ.�������H �r,�i���P5�B�כ�o�����
:(�^�`�6��LRu�V9���a\�C��_��oi����'7�0�9�gw�x�Fe8ϛ��Ė(������"�]�ӓ��[�#��Q.�"�{�,#]`t@�ͫn�Ao<��sY&��Y)0J����.�DD��lwk�d6(�Q�|��!��~����F�c��}U�vp6~�T�=mT��i�51/�v��۬���Ft=|^:�: <�^��k&��v�t�� �>�J �~Z-@_��}�L �Ǩ��������u!C\�6��(y�;r�[V&7��c4�:gm5�2��*3r�SE!�U���,F�8D/A:�9�Q���mA:$>,L�\�]F�$�
��P\זj�}k�r(�q�K(�Z^�x��׊����uz� ��͑���u[#���p�F���E�;��\��yn��IȾ7�SO���Ċ,u[	����U��z*e��vGFߦT�|����>�ѭK�!��k�u�[��p�-�x���<xkT�!�[sx��h��eG�E��H�`���pJM�5ι����y\W�㰛U2O`2���!0+�{����TW�zK�����t</@33�`x�*���a��*2�3�;ڎD;�;E()�����OML�@�&�[Dn��~>��K5�=x�}��i��B�6m�ƵSZ����F�'�BH�_��~8|x�v�'z�U(5qsk�r�V��L]�®�0�U��X��:w�n�f����e`L̎/Z���X�bU�L�*U�eyT�Y�|��$[�9�x�+Ώcr��ص�4%Z��b'���ދ�5�j����R��@�RwfX������!*�'p��S��u�.+� ��Z�ߩOS�W�x�l��y!G߳`�G�S���;|���*֌�~���u��2���;��������,���1��n6���:m����x<��sZ]Oر��U�{���uu�6��u3+8F����� �iZ�{8q�p<��s������8H>�-~81�|��\�
ҁ�\�gj��t�����4?I�Ǔ�ds�M2컉�����e�f妼���ù����_{d{u;��'"���8�{��}���w��o_�R0X߼._��ݏ�7eL%ؔ8{mG�S=#qU�T��2�����������~~<?�e�s����>?�8���?Ο�������u��L��q�uYE��^�.~}:?���t�6_�O��O2M&�����Ӆ��_��2�o���Y�A�q;\��<�����������$��������.2-�=��+N|�)1��9��:; �i����������?o/�vyy�������ڟ��w��icWx(Z	fʴ&��숗���aȊśq�@{�O�q�k�뗬���A���{�+�;��'N.�Օt�����\�s�sL�R��sO�$��� >�!.N�ܼ,p���RVd��
.��������%S����+�#]�kXB^(H=k��Y!ɣ�Vs���*;��,�"6�Z�� ��L�"A��1�,e?4j�b�.ʳR�c�y�
����5�XwkOҭu�-��=AB�G�=2��)e�C˽�u����<[�^k�kX���}~�w���䛀��nd�+�SRd���֟˫/�$/W'������_.O^�aR�c�\\-OVW[X��*O�߽��n��_m����Kl���|�sE�����*1��<�W�h���e���s��=���,8�1�/}�r�TζXV&wc�|�6�K�d8J��V��')��8,�B�W�K;_:)R�[Pl{��D�f*���Q��r�ɴ��[��u'�Y����_ �ouW[ǤKm�q��ʰ��Mwۤ���{��(�����g�'#�6�����q�?��������F�>k��[���R��b��z͐�.�W��</S�'+�.���l@�%ZRb�_)�l����<#e�w(\�b�����@�a>A�!L��Hҡm:�ݦZ�6H�hX�3��
~�\Y���Bd���"�#��c[�:v��&�P�����Ql'e~ٓ��Ȳȓ�.�K{��i�V�1β�R6{c�i���)4;�k�z�DθB��"U��������	��=6�2�A}�j=�Cv�A��\J0���L�����_:̧RF�:[�<�(�B��?��<�c�W��-�R�7�$\A��H�/����nn���ɘ��1*�1�����=Ǯ���;)+��Fy�M`|r��Su��]ѽ�"��H�������=��_׎%�g#t���r`Y�n�1�+2�WW�����(��C���択KZ��6!=o�㘷��e[����~}��'�<a��$�$�����I��OO�OS��{�����מ�x<n�W@������{YQ��DY������K��L�k(��q�<:�6yP
�u�̟3j6��,y2k�|��**�f�#���#��hvr�u��98�B�9���dO֬�V�AwC��)43j��+:R5j��JEM^T�I�}R�*Ze��q�2kwH�jO����K�n�47�5�9z�&t�Fs�'Ƽ����>5u�4W\>HM��ѭ��XR0Y(.�	���15���K�>�~�N�;�ߦl�O�O�!�;�d~������􇟥uH�kd�#���F
3��ʋ
��E_�3��T*ɘ�����9^�sb����|\�|N�윝�G��H����ZD_[KhҚ��%5-IX���Ʃ����l�%`�my��dG��T;տj^�p��T��#6�{#!�Yɀ�XM�M�e*�>�9��G}A�  #���>�s����nif���$�^.��Q��'U��>�7U=�'�[�fTq#=�dT5���-��:8_�t�r0{��SFа���۝���p`��x���;e'����aR>m��$9�lA�#��u��RF�'��bt�<�����ʲP
��랫�y���� s>��J�� w�dZO�fti/tM��Ԧ��<M�O3�3�2�3\�l����s��c��ye��ɠ�)-�Qoa:��
��A��:(FO0:���v�z3��#!5��˺eU�f#�%���5uw�:m�T��D���ĺ���k��U{�n�Ǒ�//r��ƿ�NW6���F8���`z�8x���8H$h�r��8H�$�W�~p@��J���o��pl�l��  ��멜Ѿ�|���)�����B�M�V��x.A�oɢ�6=�W�}�dE�{���1o��ԅip'G"*��#� ��)O�����EԴ�2����U�,�m��2�V��e���پ�1�d� ���
�"E�d�����gt��e��a����q},4��[�j��3���O�sZ��L��f�$�{�z��I�y�P5��w��K��R�������KjbJ���2�ze9��&܇�+	�oqc9Y�stvc�N��/��!� �=�o]6���ec��O'K���l���E��%[�ͳXw6����XŲ��f���I� ��l����`NJ��l�bF��m��;՝��&#k��Y}�G@����X���Q{�I�1g��
�k:��VT�|����sh��M�{���8w�:O��GW�t�����2ІWu	�uz��U���z�\�s~�,�FB\$�����e0%'��L`'H�Ì2u%T�WY���a�Nuw��u�}H4��@Ct� ��\���l�#УAZ��.�9-zI _2���p݋{�"{ɑ"�[���4L9a�HgP#�G�������4P�`�Q���5�69���HT������;36:���BOj�I���5P�@��]�t(̜5�~���@�F&t���p�����6��n�a`8w� $vbʀ/�2��7
�qګժ}�C��S���/ǖv��_ߵ�x���H�(�1�a��������x$6i'���"$9�r$y�!���כ��y"f�;"��L��v�K�n{aZ��,��g@�╅�ٿ�Fg$ ���/}�Gu�˳7%��M����aI�������%5ʉq�Z�0��x:Fς�5�K<� ��Wi�L��,qr��a�l�'zq�(x�RZׁQ�	�wt�n�/���I���ڱ������<,���a)��������.�{NQ��j~��U���&��.���Q���.O�H,׸������[&.W$I+7��ϛ�r�&Fꆢn�t<�������H�q�P��;?��S����/������=�}Z� �?>|��:�~}dt���@w� �/��-O�D*NV�&3��	��|YU�<:.��u�H�9).#�A�g����Q���㆝��&�v^��3/��п�k�[f�<����S,T�t����.{D4�@NI
�+,5/aXyBZO�v�K*q7��#J��heE5�C�D�Ż�,�H7�TE�eE�0�IG���r��;�7�>�������d�_��t!��NS>M.�=M>�k�3�����"���t?�כ�rJ�hq7��}݀t_� �K�*���I�}r<]�@�3��/�/-�}`ߐ�r��h8��>��]�m�&��3,`F��d.�t�L������7w�d�1���������W�l�J��_��f��#�z2W,sIj�߲���ǯ�>p�T�L7)�x�^o�.j�5�Jm%e�9�u���+���G��"�0�`Yz!Jh��$��W������9�t��n!S���}k��|��Eb$��p��U���gvZ<����o~���&<:װESq�)�ɤ�6
�%6�@(���&���@�r�J��s�Ǭ{,�=Μ��J,U{���8�eAk3=]��Dw��l�m>?\�\Gd���ã�5~�RP�rz�sV���v��u����ړ��"^��^O�a7])2��.�7}F�i�X�2Z8�,B��ݰ]�|��|��C1q1ܢb鮝7�#�AwI������|H���DRQ-�w��s��>MT/2��L������·>VW��H���� @������Aá󲔉�b�����kdt�}y���@�@�kjJ��q�3�{6�`�4�bz�sL+�U)�B�@�oج�Gе�^��*:�(s���Qw�+db2T,[�.�n�{�y7Wd� t(��C~pp��|�ޜ�z�����Cg��z8�B��e��5Α�c�\�=�у�B����X��?(���w����HO*F2'r&C�qЯ��V�/����Tw�<[�:�tr�P�;�����՝����?�77?�����#ʉy ����GH�T��]D$����Z�]x�Tb��񄌞X�n��R��^�<�E*bFjVʄ��1I�GM�*W��\�UD:�ۿ��V�����U���Mh]$�l��Ⱥ?���Մ$����ٹ��+N΀`�[�;y�w�m4|��ol�e<�[�cpa�N���{-+��sUzL���7����C����>�]z�X���o8��%z\�':}�����r4���"���΅�^F'�Z�K����?�����zyu�����������x&��uH�r�$	=�)Z������J�"�,ee���0��xJ��*��,k���
�Ws!&��h&_�]��߇t8M�c$]3�Z�~��v�N�k���u��p`�N��(�q�zTq��.�s� Ǭۊ��E�̰������ޙ_mT;k���I��9L��,(lQ?8}٤t�f�y΂�|0���r�b�dj;��o���7�3��w��oCg�ȡ��j��7L|i������<7tKD+��Zʮl��W��8[af��������[ ������@:�2�-|�^<z0N�"�E@��V�ѵp8#ɪ�����79���5�q��H,u
\Ԓ��rH�Ĺ�B6�K���cB[���`s��8Æ��[������BDIe�f@�=��2w5��������XP���|���&s�n�n�c��o�����8��/G�\�B�^o��@fd����j����6�tgN�uMg;&q�^����Y�Y���}�8��LҵE�;��C�1�G��1j�:�(|>ܻ��q�Y� �@�~�����������ׯ�{���:��*�Iw�W��^�����7��-�bQ5��Q/�,O��&�KN}r<i�]�hZH{���HL9VQ�Z4������Uq�6��%�Nw�:99���Թlt��a/oꊡ��T[��� z-��U2 t)���@��9��(6b��C�>i�<�q90ۦ�����Yt6�ѣ�[5n���,]���	�6k��Q.��}�m�.7����/q����袹GtӰ���l-2�F�18g1�u�#c%    IDAT[��]x�EQQ[�����������������������L��E2n���M�I���r:H���]oS�j����EMR�id-0cf1��	��&s�z�r��#tl��wK��V��[�9�~_�:��F^p�s��/�TW�ׯ^7����p��}~��+uM���lvEL��]ր�T�s3锔��u#
mwhV cS6�l)E��"�Fo�@P��+�:��w��SvkJ�5���"8iY�Jn�Q���+�![�x����c�ѻ���b�7,>r�k�����>pZ�B>�g�M��x�K+�.����(9^87�J�h����_����$s������'��eM���%�h_Zz��(de�g��r`���B��������ޗｃ^�fo|���_{̨r��	������K���lZʀ�5u񵷾��}���uN��g_�?~�so@O$��^��D}uc�
�A9�l:��'�zu�%�,�tS$�M�pI��9�m�ͱ���Бm���ewV�Z�`��J>��#�J�͢�>Ȇ�/��װ�h�~�� ��ޠP���?#2���f��X͋����s�� zx<0`�aQ��غ=8��?�l۲F�['~ۇ�`�]��2�6tn/j�n�t���5��i�/!�{E�L��$����C���o���?��)l:�q�������?��Λ���KNK�C�M�u�%�΁>?�������e�{V�%4���~SܨXݿ�t�m�����:����C�p�ܖ��D2���|�\"��V ��t�QM�k/�'���� ���>8����w#��A��:%YA�W9;bt�mv����r�����N0�5*C�˦�(�n���P�%っ5�d�x �/n;ŒE1��u��iF�2[�����ã���������Ǘ�~������q �����<|��V]��9U6+%$)V�7^3�Ψ�J������~=���^'���_=�&T�'��8��(_��:���������&pT���NŘu�Z#�J�8�,C,Y��������*7�	h��O�/��ŀY�
sk4�x������/�!_�pY����
��B�{£s��A,pS���_O�&~��[H1�2���GxA�q��q�|���/��5�A��	6U��&3 ��.k,���s������{��x���}��c���˛^����Y&���k\�ʕQ\��4 :�C.�\?����y�����������BNf��;��o���Ľ��U�s������E��"�b�0�UDω,W�����F��r���e�le�!��>W��M������7/�E�S�E��� ��o	�[%2z��>�Lۨ�$��q׽=����j�{�ә�g�����r��7K�¡2��D�n�� ���at̋ďd��2�*w�7���lƗ�qI�nO�Y�Alu���V/P��_��<g��ϵ�ߦ����r�/��s����>>���Ģe�L�Sɬ�xO�^;\�Y/�JٵW������KbA��Iie�	�_�C��4.\�J����]�	�ŗiM�SQ t`ȰFp×�P�eEY{Ʀ�kH��ӄ�2I\Ô\��(h�@Ķ�Zdk��a{";`iUX�N[�V������>6�Ic�|_�Go^��2�d���b��S)	�ڼ+�C+���a����Wh��Q����
�&�S\�� ���o��ޣ�Ӣ���ջ�r߻9h	F�v�N�9����#�Ǒ��զG�.��.r�sJ��-��n��n��%��IZ��������]R��d}ia�9��]g",����qUt����(J[�廉���BW\p216)�a�L�\^fH����Oc��*����h�2��ـ�uD͌L�/�����k��sF���E躴�.��q����*r�c�?2�7]N�,�+:�g�3ע��"à�&a7�|I�a8�+��u��/S`�SY�@��X0C�w���r�&�;O�w�7ݻ���D�:�;�բ��ٺ1�GYQ�{H�F���Ls��Ͻ2z�m�O��'K��6�,�9	&�r��T^j�_���љHg�h��R�ur�� �T�>�v����ư8$]s��u���g0:w��2�����dtŰ��*��(?��h�׾��GQ�Cgw��P�KG����u�{�༉'4�� �W`tHw��`p��=\Gvy����g�7�_V8`��5�w�Բ_zª�X�s��?=?����P�q�~9O/i�i���~��77_���ȳ��v3���E��kZL$%�Gg	�z���.R��`�G����艌�?QS��J���L�i�%�qIͧҙ|����£��u�rݥ�6̢%æ+���"�u12Lv�V��珗'��go���S������q'h���L���`��=:����z..��^\mq�E7I���g�&���;P�*uIj��v����\�c�Y����s�0�a@���k�������N�y��NK��C7�KK�j3��zP,�yK�v<�NŌH@�Uh�z<0�9��,H��>���\��8�6�������Uѽ������s�ҽ��ǲi}%�Φ��*���/�mJ�C������߲`�̆��\�R.;̀�:ώl��Xd�Ke1n�:��X^���R"]��_���7m4�
ٲa%�Ml����X&!P���(kn1Km�b'ݔ�tC�EZ�4�2M�E���9/i��o�)�����\�SG��bZBHO����)9�.�X���Ch^Z-�]�һJ��]��)��,]041���E�� �s��HD�O���o#��׃0��H��6�.���|�Ѭķ��v��ʮ�s�w~p0�J��������o,��].� ��aΰۘk���÷�f%��	U�F&��D���vϸ�ٚ���r�ey���^=P4AQ[�ޛ���Ǣ��1��E��`p������t��^B'3c�'�����~P����w�1s�L�?G�xH@�x��*t5.j�(�/f����cz�-y9
�(�Y�������x���u���Rzî�}���J�eW��T�DIg��y���<>��L�E?kr�ҧ�����a8���Z�l�L���]VKA�󦆼�s%�n{�w�utH�m������)��yq�e��(�/�g(�_>]���`E:�#؋����=�l�]�H ,����}1���.���0�Ǿ�8�d�]�4m��\&EX��k�EF�s��Iڙ(2���.E�C�M�sÇ�Q�P�
袸3xm�a�4z��������,k�'r�'f�6����Ձ�RL�u�;dԽZ�9���j�ċ���x"���9��L"����:a��As4�X��Z��_���e~��k���x��*��*�aU�Pw�F�|�^�Y�|0xu�#M��f(���@�__/3�H��o>�z����	�ƈ����Ή���"� �YW�@_�g;��%&�'oEC2��C�P�nE��G��EA�K�Zt��R����J��;��0 �NL�\�H~[^�~��c:�m\(־T�R.�hj���w�ʀ����hdg�!��duV��ҍ@�]����U�'J,b��i�J)>Y�b�4c���9�9^��P�S�;�<��ɸ.�k� :��W��O�]FyRω�G��"��vѯ�����w_������2k�IݓFGD���1Gc��=d@G,�*�jY��;��"jQM[98��":E_-qq!BH�!��Foa��Na�;�N0�)t�`�|:ˇ�Ŵo��*�R�q{�9ym��S�ty�i��N8�K�m����$gt�tXk>T��>�d��˻�����$ͪ�HgZ#�DԽ�D�$pϠ���o�͂fYx���`���M�����n�m$�N���u�S���f��E@Ol�Xf�#+�y�������;��6���dg��{��^4̤{��9":�m$�E�DQ1�^w������pL�}wї���~3�v����1�R4H�� ��G�Օ�Zc�Ĉ9�V�E��f&'92dSg\33̻U~Z�@���}��ڏs`��U��ՠ�<"�{��曶�b��^�ؘ̤��7jY�6$�g�Q��B$*�"[(�����Ƥ�a��2�i����g~=V��|�������������Խj�?�h$�<�k+��������#A����ʨ���۠���t^t`4�$�����~W�K#G�>�Q,��a������y����c����N�=Q����̛Y38.�����2}�Z
�]b�2�b��1:�Tܨn�6w�C�ϢYe�Lk���"����"t��i"랒�8#��%A`gH Ԃ��.D�뾟�Nf����ѶZ����b�"�t�X$�l���gX������dv�%�7���"@��D�=��H�`׺l7����������~�TG_�d�������|��Ӌ�k������������	6M������+j
OB�)0wu팀�S=�-�F?9H�/?~��\炋����mj{�/>y������F���v�7��1����K1�����5�����2�L�5�n�a�5?�K��dC�����y�R	f}8Y���$KRj2C��tb�Xᘲ�Ð��d-��J��ڧ�z���^ck��x��{�����M��������-���IjJ,��`�{<��y�!h���fL�*K�%6Tx��������I��4̤�I�b�|��	��د����fY�ۏk�FJE�/�ݹB�����8�q��@_�g;���B����m �{����19���@��]#�~�MhD�u��I�<+3�`aCv��')�D�'�L�D�*����>G���jV��O|��;Etّ�l.���ٜ�'�K�S��X,{6�8&̛3��h��4��^V����.tơa�f-K���.����:��O9~��ˉ%����9�g�n���!����d��N����1k�a�/�X1�pM@��t��{�~>�~3?�!	��Gw�0�@V/��:�zk9O��F/`U|B9�X}y���&� �i�����oy��b�`kǉzF�����+L��w'}�y&i�LY���0��~߱�iw�/I^�Aie�6Z`9���B�D�wNf��.��w$�̠��`J5p�Y�U��6�C�d%�Xr�~ՙ9�[U�#"g0�R��n�#^�%/�f{4�X��l��<0���g}��#��� ��x��
*[�
�s�ϣ �k����?zO�i���]c���G�2���N���/�?!.��p�`�q��O$1��f���?y����������QYf�� ��5�e��TX�:`B�X���XQ������Q�P�l�6	aBK����}�%ݟ�O\���+���y�� ��@_��Lݹ���'TA}Qx���\$	ufI"BD�~��܁0S�ž76U�>U�觙�{
����w5-e'F/�tn����ǻQ�� �B�@�rX8<j.U����˰M�F+��4FO��4h^5�~��[�T�����\t|I���(����Ԍ��>S�4!�;��J���0�{�W	��b�����t!��:؋��i'�$bq)B5���z*��d���g�5l�]0I�����>�s��7��l���>:�����UX��'�޷�Nv�R��*�Ʉ��/�3�IaM����녭����y.Q"��p"�j]��_��JW.��|ö���O�7?��ap�h���!�e��
��k��&ǟ��J*�T
r�jp���6�daX�ox/�zzՍ�v]w��mJ �6���!�Zr�^�$����ʇ�Nu�:��B��*����~{0�^v�.��$]�i+�B�|�v�5A��$�!Y3�80�č�����/��>�O�`�B�{}<��nb�ut���㏕|�X�`���{}���Rꮂ쮊f��<k��V����.�Yt��wy]Q���ň�����TKW0E��7\,���0F��!�j�G�Če��e7�"zf�0K���{�>����YE^����>�io.������աMǆ���}�*3�.H2��0��V����Ё���v+�u�e�#�vM��"a��:�kRn�6�G�\櫃����.9�QJ����ux�l���D�����\I
�̈́�髌w�ߞ�q}���$�k�J��j��h��"�/�3F��d1!'eUO���M�7�/BАrmN�T	͸���	e'�I�����ob~e>^bo�Jn6�F�������L�1 �u^�1xA���:�2qH���|�",�vfX۞5��ը���t��%Ecf���e����^�	OD('VTJM��d�� m1�d���Lc{6�=z;��{��*/�f�lnǚqt�:��!��E����G3����o��M�>�<�R?K���[
�(ٙd\j.K@�����]�����K�B:�ρ��q%A�<���Wf��<��9���x.��tap�e\w.�86�5N���|\�����ʗcH';]'�flq�vY����R�X�ɔ)hW )�>�p2��������,h~hi�����Š�؞ւZ�`ٞ­LUt!U�����ё � �����jtf�jiT�;!��}��+��Z��1��fA'�юw�ƌ������A��	\��E*[De}��ͻ���&�uݘ��W1J3L�=<<�O��
��S�4��&�g�k
�d��ທ��0N������8��u���R!-S�����<@e��x(�E�Ǖ�ά��ڏQ掙��g�n�,�q�/���n���~w��S���9E�J�%]���um���)�Ƒ��j�^���n����:,72ӳ�_g{8�T!�\���Z#3f\5�5mƒ�bp[�Yh����Z�Y�M�����y	C-1�c�HI�K�� 29{ʳ������Ε$������/��?M����<���}./���@����2t&�L/�a�l��5I��E�8�x^�kj� s�E�u�	���
�	M1w��=���ipM��;���>6ʵ���]�m�g���L�)��%&<A��	ʒ��ݏA�ھ�T�cu=���QM�SZ�T�ەJ�Vi������ui҅6�'��uN�xI���&1G���&}�s-�Ȱ�����W���=h�ӫa3������;��{��,R��b�g�T��7���9l�����>�x�M�D���_���L1n�9�᧔������tF��j�W��-P`WTl�$�/�s}m��� ����qtN+���PO��D3c{�MPv �c_�øi���Q?#D�o��{��a��+�9^�)R�˖,Rh{��Y�7���ٙ����_^^�F����vL���ϖU<���������Ee����d��@�5��=F�E�V~׾`�ڠw}y]�p�Ei;V���� +���������0�~�Cnε`�k�=�/p&�[x,�.��667SO4�峣�O�_)���H3(�����	��o���`�%s��y�s��PE^P%l�Q�~J5��� .���t5�f��	/����O��2�N���ʸ����<�Y8��^�t�?G3Nd:R|���b
3hҳ����R��m�4�a��i>��'�z��-�^�R�_�<l�)��{Aρ߹o�����8k�7�����aǰ�1�پ�	}����f/+��t�"k�Λw�0fJt����;�6V�׿|�����/G�_A�[N�o<��C������ё��JJrD������ɿW��	�o�����Ғ*����/�n�d�X�="SbL@��Uz�t������f�����w:m.K���}Ӳl�C���.�#E�qb�Cmg�p�d���@/����P�t)���vX�M?�V����uNHJ�~���S��k��c�j{�F��,[~����5!�4uV��8$���Ȕк4QU4��2Et�`�,�l);�������{�}���| N@���Sp;8T�<�ܷs16��$�$J�+X���B%�� �7`�cϜ{n߫�`fؗ�*�����t��j�3�3�/�ȿ<��g֊C�j���еU�& �����m�˰��*�����j��f))�v-K[ }��hѕ��z�]:���<"ZΩ����*L���Ϝ^:]O;    IDAT�d)��J�g��A�[ ���2���B�G^�������O{J�BpO5M���8�����`�joea�ć�]���(�Aӂ����}�p��B5s���l���f��{%���LK�;E�x�'�m�Z"oq���l}�"V�no�����c�#��>%�|��0������;��вz������lc�5GRhb�d��WK��݁��¢/�-:�*�)�t��=��BD��lʪ������$� ��� .@JBTx�[՘����q���QwrL�Qe�%�M-�px>#��6� Y!���4ɂ�<�)��h�N��G@���z���"UQ�I-�{�y���"�]-�}X{zY�z]#���c��4���@�h�	#�VfY��������������������1��_�H<%��>� ��E��]��5G�_�:����Q?�'�}�+j�aHd|�1K�M4�Z
�W���	�� ���V&膺҄{O"�?��u<L�M��נ���G�H�Wj��DD�ɟ^����㊹|r�/��4e�� ���4C���D��	7�$��)$����9l$� qi�:f�м0�Nj�ȣ礷�W��GG]�Θŗ�2����y�}VW�X�~p��,1aKrv��tF>zc�*��F�}�����1\�����>�kW=½af���	�f�ڼ�O�+0�����$!�췘C�4�߄�&�GA����S��D>�n����q�ڬ���kaO8p�-A����xr0"5�L�q��^ԡY�3�孓fN�>���}�Ёj��v��ẇ�AE�'dRR��n�sё^2E�jf�W�BmxV��\~pg�׾mk���Qg1{��(��o��ww��N�ܶ;}��	t݁��kՉ�7��,t\A���eٸ�u�wӽ��r���̊GB�.�f�V6�@U�''�մ; �n!���&��;Dݹ�.Z�؀�����D��?��i�E�(��ƐtK�<�W�,<����oG�=�G����`���=`�_�K�"�zN�l�Z�]�Q'2f߯��e�eͳ뢕5{�ϓOD�O��Įa��mX������m �u}��J�q�`��;䢓E�#�m�_�\����CJjS��@s zE�u�@���"�!!zr�G鍈�+��*ɘ�VG�B&���^f��p֓Sw�1�@�����	�yW�ɿP �����y�)�--
og�sKAl�q�c�7���Jn���;��`�˳l:�Zf�W�Yx�,`M�'�Q��D�,����pZw,��B���z�0�"�߶x"�"�X󌺯�W%����g�qjQ�I�L�5/�ݛ��q�ƹ*�f��DQ���;"_� S+�q0�Bם�N7��c;c��c��P ��|���gEď_yp�Lj�	�{_��9J9��T��V�A�&��\��{�؏`�O����yP������$���>5��Ӄk��Nv��fu3k��,LW.߆��x�Zu��iޢC�.$�8��Z?��޼�w�X���-���;]� p��}���8E�6LfRY˕�w��Y0��F�dOW�$;��<�*�Zm<�XtLR5�(�Jq�l�V�u���@=
����YgF|��g�1��!�'�j�eIQ$��;ݭ������A�l۸����e�}�[s0�_,�2]3Gw�͟�_��֝�Kͨ�0�'����~����^�M�O��7��5GҬ���4˶����y�`�nw�k�5G�N��a8VGDݛ��N��䒦�����,j?���'Q��>w��~��Gt"N�J|�{q\�=:z�<����*-��t�X���b�b���V��?��8��ⷎ���%�h��{A���9{�~�Ry��awtXr1beq����L���;�݃J�n�!F�����`a���ڊv�n��uEwd�*-U��~�<������~+?�t���{�`�g�=����<Ƀ䐚w �n8�3Ժ�H&�l��Y�~�57���G'��M-�ã^� �%�t�)��#�Qw�Wr��\��c��w�q<f���8���%�y:��*uCUQp'o�+5��p?=�}��1����t�1�XOhV��>m?�ɪF�\�!��Pi�?��P#3�6�8��8h�c2���l�D]�7�E���a���?�.&88���X��O�{���zt{|��շǻg/>���og,�<�k(E�,���Q�Zm�-d׶-ki�/��V�d[�����>�݂!7a}�[��z��;�i��O��]M�~��OÐ�t�;�O�Ӵ?m��0���������OQ>_T�CGv�Q�_V���!�k���Ӵ����#�U�>�ҝ��i����c:����A�MV���%C%��R���/�Aw:����\N�,���]��� �t��2�����2��C���k}[q�T� ؝|�������﴾�ח/��֟��ǟ�c�ZZ[׵0�B��x`��=0T�d�Ih��$��(��ɠҴ�Ji9�S�nw�r�����)��'t�?d�Zv������~ӿX������1��,>�5@Zpb��"�ޯ2cU��؏~�/�-����U�}�|�2�-�y!?X��v׋h/��e�\��X-��x1J�+V���xZn��4֓�X����Qq�j���}6��K\�$S6��bdr1�����soG���� R��!�!���Ys1}��.��?ǽ1]�ٛ��{�����w1�)�{�8��{���m��]�>�Q`Ô�Գ�����9ڝ{�����'��O'Oӧ�	ʓ�����d2y����d:�k~s��"Q6�Q'�9Pt�+?�@76R���@?җѦ͏q������'/P�!��@��4�)L�29?^~������������寺Y��^/�A�j?^��aTT�������m_�y%6��g��_f{����3D]�����]N��^kQ��z:�P��l��g#������r�5���y�>�~9�����o�������z��Ö�g����>�>?�rw����3�_�o�Ǚ�Yjw���amjZ���{�JU����~��z��6&5��N:4z�t}��	�L2��}�'S(�S*����1=�-�z;�mI��m�\]෺ M'��nVx;��B�����e5�kp�j��X}C���n���f�}[�b_�x����j���t+���*��i�2s��d;ڎF���t4��3�~;�g��1�G�n��L���ў8=Uy��Ў���dq6��~��~}&�oP8��c���^�xa@����{��L��<�`i�4�7��ٻ��8)uQ�я�@?��(�U}sv���@pti"����Be��ݽ��5�a=r���:�vV�T�Ў �塋����/��[����G�T����������������=�{��^֬�����m��b�r�33a�y>�A�K�����&�G���a��I�-! B�(�F�o#V�mG��كD��|`2s�|�y����������l>�Yl替6s
77l��͏�|�c���f�؀��Ŧ_����Ǒ��;���V�����%+��I���#}�O,q��"^o�ج���P��F$Q�U�]Ҡ��6M���.�<�*��h����J~�e(�\��)a�{"4i�ēg���W=ʱ�_���Ty�H),�@��H���2^��� �8������Ϲ�[�q~i8#����0ъ3U�I)ն��m)d K�vk�^�]Y��eU���j�ۭ׻��n��xرFv2]�>��}Hp4�]���*+B�)�_ݏ��@o'��E���??�|tc�&F�	\`�����N��I�$m�MԎd��I[��(
�F���5m �ID� �R�X5Qg�2>p��)Σ�pR�F[�I�%/��.��7�g���
ϑ�
�;f����MA4��ݴZ�&��a�՜ĝ.�Db�w#ʌ&�U��$�#�sa���U#��}��8>�ĝNV�8�q'>�:�<;�d�YcaE�V���1q�CtS�?�u?���L��h������4:�wk;���?}���#v
�iJ8�R���	si��y%r���TV�@o	�V�%��jq���������Zޔ {P�	\� (�9�5R9}6���r,�P`pr�T�fn#~0��-�E���C��ƕE���x��YgM^����R���:�`�
�m?97�^��88�0���1m>��ͭ�m�,�e�qX�4�PߒP�w�
v����HR��O�2�u� ʹ�!s��׎�ut�/����Wa �ᵄ����o��DT�P�$��
����=��2�1 �O��VA���Q!u��hI�)(啶��9��b�U��t�����`���`,(�!W���8��%�3*N(M('�)h�l$#�'сQ.���ɂ��HE'Z$~�8;�`��������%����~��C�e�HF���֦��sX�	�wL�O�!���／����F?��i��S�@/u�|��K��ӌ:!��4CEr�7S��� C,
���H��N��HNs�^
��H����J�0��K*u �/�cYK'�;� &&4<��j�?,~��M6��adY��44��
�=�X�Ps�
�,��+�&5�C�H����>��(`��.h��:�#��($���˸����yNZ��P���H<�$9�J��6����>T�״*|��#Џ�e�oK�j�Ǐc��/Y�2\\�HMĨa6�HӒ�D�0�x�%]x(b�T*�`Lp� $ Ex��Ō�q�ǏD�o�LP�RX����p�Ch����\��U�^�V�(�>(�
�������da�����Ґ��K	�Iqq���;�%���c7��[��n�]���!��~ߑӲ�@�<֏�HV��|�9sFI�У���~&�s.r���� 1�≩h�������Z.��)�7�lܝ�q�4p�̸���
���
�+\�zm��ē���5���VN�D��vy��π*9��Q-��oS^�F7��m�Uv��3��ZM��l��"Gy�	����;��$�n���0�)�L����
�`��	8
�G�6���Dƭ�t�ߣ���>ŉm��	�ao�ueJ� �1���x�zE���o�b\l��ҒeJ�i�^���`��Y#�R-�=�E�f�o;0J�P�ؖ����ak�8kA���	�|�`�	.�΄0�P�o�z���������r6��њ~u�^`��m;�o<
C���&^ʆ�7��3���Ӫ�Pu��Q[\��2�:Ё�W]�{ ܸ!@�&!"�s@���i��Lnнn�ډ����[S�.3��������:�?DE�"b����x,��9��0��/z��4���.�MI�����C���"O�t��څ�+�?�dȹ��8]�7�YHÜ5�0M����ot��z���S��NY]ߌ^۔+�mZ�|���V�6d���2=�#:YS<W�{V�~E�J��5^e��6�r���Ib��q�D�Q��w؁�Mߝ����v���P�hnF��ı�(�Nˤ�ٯ�n�b/���6{𩐛*�\q8VͿ��cXd^�q\i���BO�g���1�>~���1B覲�e>&>t�ew��I��8��f�y�6���fK%I̲y�TR�vNsV{��Mwݘ�wX�0-���(�Q��]�U\��dB�ZS�ub�!C[�z�G�!���9��	��L=k|�̰�����ւ�-x^YT�ȷ�l�]�$5�$Q:@Eʀ穀KnY����	؛*;W�"m<zЈc]q���q�P�%p>.
A�֡�G�~_�v��P��ώ�5�eN�U��ĉU���{��@����t�#6��?@籿y�6��l�]K�=d����>O��0�}z��;��u�M�5���>3��#�� ��z�oqkX��8VqҬ����x+�T�T�Mׇ�Po�QS:ƨ! �ڍ��\�P{���P�(���Jr�Ǚ���Ўo8����Nʤ����M��B6Ѡ.��������$w���
 �>&ًNG��/mJv�뒋)����ȕ
�����jvT��J��U�j���0N��s�=�3�(�%մ��oS^Lu���	���o��k4rC� �wu�fY�^�շ&��:P�'�m;�1���5�z\�moכ�z�6K���ǋcp�#S�a=m��QkKc^���і��]�be8���nWѷ)�Z	¥nz�A��GVW1j�ZZ��k�F~d�V������j=1)��J��L~|�����}�)�~�U���#��; ��B�ZN�;Tw�JJ ]� }S^��k$��*��{d��i	�ܕ灃w��ǩ�<�9�;���;�����nPX�nn�~�֛j0��1Gv����ټ��$��?���{���yv�����Wf�G�ϸ9�����9��jl�B/o��N[#�i�JO���,��n���˧���b�4����r<?��v���O8����y-K����t.z���4����nǷ���v>�_q{���|<���WU}.�.��$��\���v>T�v�I,�)a�����)/h���2?�Z��+ΪI	�p�΃���Go:�ѨS�K��*p���-�hŹѲ[����U�o��y�<б����i��=ǽ����C��G{GG�2+���la9<�CC﨏��=<��m�@z���}��)����;z�v5��-;�����Vg9z���G-�/_u���w:�W����I+>�4J�J��n�ŏ��\u�V������U��}���W+6��oWg]Y&[���n�f�L�*�{#pw��Fo1���ne����)/��ۦd�TX�s��s�eb�6�[":6NgF;��AU��N��M���O��X��y��/�@G0������<O��[5~pк�q��;�M����AU��[������\��ߝ���,��/�Zp�N�����T�I���`}�ܴ�d��`���e���n�R��{oZ���|}?n>��}����Q��{�q`G�H�x�׻yO�d6�ҏ���)/�K�b�VN��~k��%�W	ڱQ*�X|h�>�-��pu2,V'�d2��b�_��U��py�+x~9.��~����j0-��X��Ħ�(��{�vNzSFIڨ�a����,'��z#&��I�)���0�Tb���Y�n��;>I|�����8�3}ԏ��-���������Fˢ譊b�Ϫ�����|��^1L���w�ܦ��s�q0V��W��`r��d�A�g��>����%Ǫ��6�E{�K.�c�'Oٽ��7��@��*�D�m��9�2�s�ϵ��L%=gt��t��	���h�����ò�m�~����:M��HD��l��w�s��Y��@�M��w���_�<<p�������������+k_Y��������]1�$��޵5��]�aLz�L!��ґ�g�%��)��	�%V�1��r��`�&��=�8��IM���_w}K�=}9/~b��Bb������ׇy<F#���+ox3�ә����t9����;z�ca4�C�G�D����߼J_���Ǡ3_ּ�yv�����k�>&��f��Yw6�&���u0�� ��o��ݫt��O�Q�r�8<�id�7���߫T��_�V��Z-��)#�����.�U	a�
�hшz�{ϫܹ��}��ٹ��W@�꺴�n��{����w:���MZ���\���:�B'��̨���q�fZ���r����Ȥ�U]�� #/L/2��px������oo߁����m��"t<j<-z��W�]������[|`^�w1���_Q��xL�D�C�6/���qO����ʢ��cFݑ8�He��3�'uD��p�xP��m���7캮m����3;�������h�4���d1�{@�ܯ����	Y�xH��"�5��y�v��~)���K,� n�n�
�5n�|-�B����tZi�U;�����z�U�\���P�>������ơ�B����k�ܱ3p݊׭LU�+����B��h�%�*    IDAT��u��ó�������� ����MX5�L�g����zd92v���Wy��#�cRV�ZV�1�^7�������';�H���Qc]K���}�Ң$��(+��&Mu��$��i��iɶ!l�d�^�U�EF�@x-��]+�u���Xi}	�V�iJ�O�#h���;$��vk�;d�#z&E�w/��3z�0�qV���E'i�M�i7�p�ˤ	*j�n����BC���7R��W�����z:fti8��l}��t��+��˶�]�x��T����	ǥH$"E���!�p��l�TUV�}��]A!�����ϋ���e��)�
��ͦd�?�ݹ@9ˉ��:!9Aww��b�Xo��b����	��ѳ�*ƍp�]T2��̓���p��*͗ҥ4��Ҋ$D�K�_˦%�:��/�v����zR�]w|;+���g�
:7:g���#6�����~�����<RV�<%Oe*���K׷���S�ղD2�^j���|�E�����4Z��闍�f� >z^p>�XU�Y�Gl��ap�#���~�c<w(Ѣq�X���d��-��-��$9��;I<����*N�:���X����KD����y����f2�l_4��)e��d��d�%�ظ�i�v����׿�!#g&����]o�pX�b�S�A����i�����6C.��~k��^9&�:1�&�7/'׮~�ka>����7�m&�T�S$����+��b���x\F��"v~���qBB�������h�S^��!�^����|K2��������7��DYt6�>�6�^���|��/1^�tGz��j�`�q�L�!�{xv�me�B��<:ʲb�&d�Ӏ��4���2Q�$�>�>k�����>�#�CCe��?�N2׋1� &��0�0�v#� ��R"}֭n y��"ŷF��p�{+����K�k�i�n/7�hC��J��|8���+L�Ƞp�"R��!�8]F��u_�G�?�Qa�\U9���^fè�W^�j8%�> ��w�(5��:,���yFA q��b�~�Naё��ɲ����vm�w�c6�cPCh��Mf��]*m�����41y��Y���G�w�r��ؐO.��/���±����G�2L�A=��[~d���O��P�yLZܯ�z�br8w�D����������{ �j�L�����QlKH�'��pHR"[k̓��y����j\Y�~��X��Fli��`\����b��Z4���QE�o8�}st��Dׁ��L�M�kF���%!���b�8M�G���\?i_��8��ur�ҁ�d��Xz����l:Y*!�*Ѵ���~������!f@�D���4C=�Lv����b��c	���v'eZ�On"�D�O']�XZt��Y��kZ���@��a���W��=���O�E?��?�5�K�K���..����w)���OY}�Ϣ�FD���Y�$P�!�"Dݻ�i�ε�n���4�0nں�p4ny,�=�/Fd
@��\J��C�Q�����<y�`3�L?!x���g9G��"X�$y�L�`�i2��Η�W��˘0��"!����M t�a'��?N��Yb���<��r�ړ��jLH<�������{�p\���B��hмހ6�n���0���.�v���l���DM�j!�֛{ū��+r�:Q����o����W�G�$���\��t��A�u�a$3�����lbB7a<��e��qۓ��3]f���r�����A}�Q?9l��w�G�T'۝KZ�O[��R�(z��JOKI��7r�]��u��ߟ�tUD�2�"���"|�]]/��8��ԙ��	�ux�����D>�F{��N�f��ز*��zӟ���xIL���Vc������^�L�1���}�+JU'P_&�F`�3u�г�
�n�U{4��?pœ�P?��X�U.!���B[�M�m-VG�;�f��z��#��\g������MD�|�����>|�<�qi~uI��}P�{Dғ�5/�����>��f�aa��� �˯Eܑ����J	je�qТ��u�`�m}��4*T����{n���D���629�9���܇М��ы���������Rt:5mc</�}�Y,V~y_;�)�1&Bȣ7w���|t'���(���uH���}��v���{}:�����71:Kw��!R��郁>2���o�&��G�����G��|�<��8E�|�����?���-��
��or���!S��k�6ՕʷW�cK1�EC�����k(7��`���f���	W�����䁙\�f����PA�2&����U��'j�E0�����S"Er}�$}�����Տ��D4��5�=<�s%��<z�L��[�Sq¥K�>�Q�3ODs���0%�)�M�C[ �/0��"���#x����*�7� �2<��Hs�a�fעO���@�	�¡O?�*�!y���<hz�<�ʃ!x�#(���7��B��H��d8��zQ�ӃGD&龲���+�a��zL�SU3��=s���egn;^�KW��8N�coKw��u�7�	26���.�ET��S�(��S���bZ%��n_|����7�|�r����f[��5;,$ݳo��Ok�ݲ#��)1�	�'m�n���+��b�!�G�p��q?l�$�n�u���/�s�,�^��B���'!��[ ��˲�#� ׮�^x�������lYC*19*<������Z�Ot��`|��M�z�P�GA�\�,���f¢'H�+��$��0:39�91�8䪐$� �"�s,���p}t;+:Q����Q�=z*5�R���.�Rj+�N��ײ��ս����Z���=���%���%�PK�� :1���ƬH˜9=����u1�)\x�yL稠�4NɡJ�Љ��XA6������A�;���u�~Ÿ=�v�3���f���Zk@�n�+��=0���Y��ˣ"=>Arbo.������!��+����7�^��*�<�&F�	3�$�D�N�>�$(e7z��^�i_�"JP��ۺ��;�������N�~��X`+j�&�;t�@T�~?R2�Ix���۹��?���Z�V���}�NG��[)"~��1��7��qg�-�8ꡣ��N��k��M����V��е��)�~ A>�T��G[��N�[���!�-��f�w�Ǐ<v�
�1���w7��]�f���7F:����=��٣��X��5��=1'1�ʛӌ IBX"_4��zIF�dl�ȣ/у�m�����_��NӼ��o\W��� dԉ&�,�6v��l�ё�g��ߎh5��4Iw|�hk�m��v4Eޛ~�%u9U��v����|��<�>��ս��vZ�F�ƶҏ��ŭO��B��sH�SXCG�;7���$m��>�:�zd��u�^��p��\h��N��>�#�|s7y0����t���ܮw��;�n胑� V7��鞌�����{s��(���)~!���{q��(�����O����28 8s}����l�)��%ㄢЧ���p�
���S���lI(���fX#|q3Ar��{o�w�.���$Xnm�U����R[ȴ��?����y;��]�k�j5{՞N������K�����ۍ�o��r�"u|2y�N�ԍqM�é�� �����և�Q�`���دr2�]��m��`�|�7f������y2�Fo��q��C�|�A+\��c���Z�l�a������)�e��>s���]Z�^�O}r�$ЉE	@G2�ͯ�D�����<�3s����	�H�+I��!�����4bv�a���J�XS�0�4�V�i]�H�K�Ɯ;k$��ܔ��F[�����''���"W��o�g[���J%���to��qI2���2�%���-p!�Ю���1jXC ��d6��A`}ty.��G`c�Κ"�|J��?�h�ѭ;�J�\�K���A�,h��@}����}����!�Řke�=�vAQ,�K�O�:Iw*,BGٛ����5I��h�(��B���3G\u��,��W�Fw�B������H�{l�WdJ�ov:���S�S�«˭���tGw<�Y�2p��d�+��\:M$���j��G;=�(E饳*-	���nq��k���ef�C�c�60�{ohi���-�5�nQ�����rޗn'��MN�q(�t��%��>����cZ���NH��D�&� [���}@? �KA���<�սq���-�����O�:;x��K+��yeA�=�c\�����w{t�S����n�5n�A��x��;�G`ώ���qA��lN��ee�<�c:WʕԒ?5�J�����U�&�\4�&�۟�{��Jn1�j�����/���b�r���t��T>M
���49�n���p1wR#<-k@Z�߸5�E�?_�<�b�t��q!&	O'.cs��w�u���Wl�n��a�ɕ.{v��f����;�t�ڔ�<��e���^�����t�C
����or�нc��k�uG1�u��t9]����c����q8(���'��	]\���'�:88���hM��ȣ�p{m��Z˭�?����b�V�͞#�K��s9����瓄�.�۩��2Iwd�˿^<��8�\
�>;�����hd�h��0���]mO��L.����ρTP��VEi0����6-̱�����@������~F�x &�	"�5{���^�Sm
F��^6���G!qfV��F��Y��j��ctM��n��n�<��t�?d2y�o���Yv�m����lb�c��iL�"�{}<�>v����W|Z. }p���QjNU����V�Rb���*!?R�R�@9_��J��[�U�wE��@���PnX�<�N���Wsy<�����@�B\�x�D`>���.�(s߻���e&3�K{KwW:zotO��L���V����J݉�w��5���H)����c���������i�r�?�s.<�R�o�C)ޏ�⸜�"�Ω��1�<�":8��9����^7l2�&xgzj�;�F�?���k�}���������)���o|ڟ }p�u��xHGO@7�|�UU���D��=�#�,G� C�z�j�=�o��t����w	�n���=�ȫ��nU[y�j��54��u:��\0yuG����\2O){O�"�g?}H��zf>-���7�V)�c'�;�J>�Q�k��i��4��� *�ηjU�V�Z�Xl}���8+u���� J��hZœT.$mp���2�|�b{�����cp{���Iw8{�I�����6����ر���!7K�}S���Db�Џ��Q_���؀�N9:]�
���Y��������<X:��<����Ky(`�e��RG(m�M&!���Z�2^�&�:d��T��k5�/ގ�i��S\���(�'.�1��YO׃�x L��e�(��댞	$�n���{�tfs��w���SD?Y�i*��cT&����V������(�ն7l�^�f6nG��MDN�Δ;����4g�9�>u�ʸ���!�ޱ��N��=g��B~� �9�(����c��alqw�>/eH�	��[����� }p����b�hek!�r�d%�hn���r���"��l���.�Yc�K���_X����bi���U4���&"zS|�����^m����)��&	�`:�{P|�����t�Fr���>��ո�L&���N�~�|u��Z\�!���Jh����i��a3�^���dʂ��l��F�܃uk��q�a ����T��؜�ыџ��)��TU�|��;�G�-�<�Z�ۯj�k��w��|�
�C���t��a.S@�~��)l'���*������ŨK�*D~UEN�b�eU��'��6�]}�k�g�E@�`Y��h	���F���y��]�`F���fV+����ԃ�� %�=����ѷ���	]�'�.�_�(�g2D�7Y�N�_�������z�5��ëz��8�Z�i]	�8�b�.�?P�A�r�#ѡ����k��E.E���s�������aF��ݜM ��\��]z�@���1���ڍ�F�p�u�0������<���_�>0%��� �N���7$�Z�$�/��5���nh�@�O���c(>�#�q�n	�!��xXk<���rc9+測qDopꎊ=��VWK7��s8�I����q�f���u}"��b�����I8��H����dW�_�n7680��_H�����P����A��m�1	�lhy;�ñ���:�[�x2ƞq<�
��~&
��.�������z�!u����
��=�"�;Rg�)a�>E�=k��CJ�~.��Q|߹� ��?�K��%���{����"<��u�E����q���	��}K��|��uJb�<"+���^���Cpm���2�Zv`���`����`���.���Q�������=�BR�^��]����*�Tǽ�Ct�?Q��N$nQu��Uv��n�ݵ�y\7!.��:�,Gb�vtC�1vS��M��K��~�Wݫ(D`Н"z�Ȳ�ڱΎR�V�!��T�"���TU�\fQu�VKptz���ǈ�ay��p��`|jyHG5��mhR�_+ފN��a�W�Gg����a�����.�F��Xv:+{W���g��/���0��0t��W*<��&���yL&>��'2s׻����UR�'�Y�"�N�;�!9��7.�Kzƭ�����b:8�����^s��<�W�U�>�}U�G��Cـ�=�T�˶�.�0õ
�`K}n����t�Zw������G*O�1u��:�5���	:L =�ǣ�]�2��.Qu�+��5z�@����ؽ���u��ux��BI�y`	�篧EN�ew���D\d7����	J_�o��+�d{�n
:�X6��.�V�_���{����s�I����d2s�)[�k�����@:	�sD���p�A�.����難1+Q��h%���8��I��]�Cö,��X�h�M#�d���s С�����j��<<&�N�;��quo��kfL���o �B�XZ�H#J���o�)pkn��GO�v��ӋHݷn�
��a%V@��=uռ�(zT��K���r��^-���R�����P���O�e��r�����2��=�,ؙG�R���/s�x�26��X�g�ub������z2>�����kI����:v0rD?���L@��ހ%3�,����Am��|�������j�ʺ���G~A7���9��
��k�Y9��\�E�ʸ��#��p��ca�Lk䎇X�>����1������=�1��I�Sa�)�A�>8�;_�94{(�L��ZH���`����u�Q�B1�t�3���HcFl�x�&�ܡ�����݆Є:��l������R Q����������| �I]�����'��)H���k�I#��!��٘|��L3\ҭm -�j��Z���ب���*(�e�.���?�;�y�?�K�MK��̙s{.R��.�}�MgAH_�#a�~{Q��.���+�9=�e>�@j��4a���+��}J��~�iu��ϝ�9-�ǻc���Nw=��8��Ӥ���[[Q��.���kc��'`cP�G��sd����уԮ(�1 �Q�]�%Cu����˻��3���A�,��Lj�}��jH��
gQ=|�����+�������z�vN�������c�4�5��򺤱�b@�Xa�|�!�Gx�d'��ѯ�����''�G�x�~��}�2;+/g�kg/+�����[��W;��{�7^Rɱ����O��K�����n����(�5�g�N���i#S���s�b�nC��`�Q���Cr��\�M���S�F���S3H=�y�X� ���y�;�:�cy��Zz��km�KuERy�.�qԣW >@��ѣXȝw䌂-Ѝ���f�N��lq���ą�a�4��א�)�A�E����(ݳ�d�Ŧ�k�X���� �gGӏO��re���u��:8T��j�if\xޚF�j�    IDAT:�A׽��ₙ[��.�"�=��1�6̰����Y��j"��x��~̚qBt""�2�Go��j26���x|�II����O����!���琒�T0V ��+ݽ3��>�z�jId��ԣk ��Ak�=�ҝz�A	�V,�!��"2�������ѩ���g�3:�\�F�4��NO�qb�����R�y�'���}/
z:�wU�R�ß0g��J�^�(�)�K�4��C��q�ű��B8Q@���P��v� �^��#E��|t,��f����Z�)5��l��_|tw�V�E��1�6��G���s���tL@�����d���ø͌BWL=��Z^���zم��q+���T^���G�2�ۻ�v/K����B-�y�;�d����Of�w8J�Y{�]������ ̼i�<�2+-Y�&'��l:}t�[,���x�����Ź3����!'�,��=e�{fޯ��(��^�S�{�ƻ����	����M	"�	!	�da�Z[��zM�_��ρ�cd���f�<��0���u��r��Σ��O�	�dX2aӠ8YQ���N��61*.o��7���θ=�7��o�[.��H�c� �Hjf��KNn�c�^�1E�$�a0w��0��8���f��?�8�2:��k��y�㜀��iz}{�I8/U2#���N���J1tzpNG��m�iW�2�~Lȩ��SKǹwjA\rp�Ŕn8Ї=*�M,՘Xg'\��H� �jk73�GcwC~�6�Sq����L���&�4D�;����'��<��\b�5�i��j�O����V����S�����]�f\��\jfw�C��(�}>VE�n�jE0��N
e*s<�e:����X8
R@`��a&�~Z�v@�a��B�����`�>���6�Gk��G�����Gd�,�q�v�{���>���YT `�<�N����X��0	O�K
��0Tܜ�����3:zt��}uB��ݭ��BIø�N�w�e��T�P�SEC����s��8�U���{V% S}$��ģ͹T*�ҝU�4���w�yg\ø$׵ ���R��,%]�bew*J��Zw�`ʗ�Qn���es�n���O��lD
���5�u�Y8�k�8���ѩrN	=	bZ4����]������iu���1���#+xk{{�-�q�/.�&�^�P�7�����a�E��A���Qځ(,D�L��͑>�M�}*�y����Kvz�f��pWu~/�{�V��^��8o��م�fX.��5�c�u�_C~�˳������ji^��1�byK,u�r�s��CT�OH��� �D�������LD3k;`��d5���W��tN`b��7X2�k�yk
�6��pf����l��$����j�|]�������u�w8`Wg��z]���+wAMRe��%�Q��f\��rzB�X�
�ayƚ��N�~�U�-�Z����/5�dd��O�l������}�P�����ߐ�i�Ȇ9�uC��YxB��M�����
��B���%��;c� �s2��S��ff^���iTa�\}}�S�v8m���7���f��q�� ��ڴ��2e�f�)���_��f�=:�@?E���zZ�Cz��r}]�V��v����h�����(�OW�gv�}>��?v]t{�Q�#6
��&���90?а�	۽?:�����c1 �i�b��ZS��"Bԝ�����K�K�ǯ�{}21�ƌ��q`���	f������c��)�_m�+���^���2�F�9�kBaf1���2��>��:MS�����Kp9a�5#��J�@���L$2RX2Ωa�fH�J�_�(��N�������9�1b=M>Kc������
��������ٴk�
�X�����uB��]2��]����@$��w�r��v�r��Vm��.��|L������o��M�ٜ��X�Q���v�ӿ�;����h��Խ���=b����y3w���ꖥ+�1��;c�ѧ�K��9�:��X���>�q
����"�q.��#;%D7�Y!��4��5î
e��S���A�ˊ��=�9��<dK�yږ^�M_\����_βkb.τ.��]�g��ջ+.K��59�ĭ��'͎X����tu�/��	����#��0r����3�<����۝�V���M�?�l��*5�~36��s��/`���?b;��2H���=�\9�B�NY> �5/�{g|��+�-ޣ�.�1]G�K��"�0���d��'���d��A�.&�A�҇"�O�>-�7�������7m,�2�E#��c��-�&eY-фKChh�Y��)a!i�3!l�U���d�L�T���=�{l�|���'�cc���y��;��D�� �m��:�������뛛�7�h���	�!�=�Wͽ�|YH�I#�i������8\��K<@`��N.�\��z��Iߡ�8�c1Cӷ/Vg���sɎz=�z�*=�r+����j�y�*X`�8���9�v��t]�rt#%�Dcy@7P���F'O�9��^cL�C}�ԩ姝"��)M�,� J�����5<{d�U_����A]PQ�"�3�
�5$�1i�	���- ���{�)��<�i��FaG��L��vU=�V�3/�ʝ?�f�{�am��3B�
e��u*j��y���h�^^9����g4t�Ah�97��-��	����{�'�k���Q8 L�PJ(ji�tM�U�0����/�Tݩ>�Ef��qU���h��?���s�b����p6g�
�R�k�VPKbR����~Ā~��d6k(�hHJ�I���u'lCG�T��� ���QK��$=�0�)�_yvU�;\�R����lt�C��q~&일Ŝt��V�L8��~ǀ��!��&Z;%+ݳ��p;�(-��£i���ߡ�:��FL�d��ˆ,l�s�'�Z`�=Kz�h�5MK���E��.i� K���KR�]b����x�*���o�?�N� ѿ���N���H����`�A�
(�I��Jf���`P`����7ph\5��MYɇ����xf\�W�C���P�΄�<�h�_ۇh�,Sү�%J�� e��%���7��������6��y���3���j\I���`����"��U�D�_4�&�M��sg3!��EJ�|�V������@G���o�`�i��ǚs$SQ�}�0)1AU���A���7�=�N��!�F�4Ș�b>[����:�\5;�+�!*�Q��Ͽ?�Mϩz� �|� �<5v�\˄p���M��`���ٴ�z��^`��BaX�
�b�n.$�0�@�)��x�����d��J�Y6R?D�_4�f�k1�=3��L՝�k"�ΞNrC�Z��!�0�a���-T
���3b�4��D%�^�ב�-���^�n�a��uR��\6��qj��k��f-m�2]/'��F�y=�|���ZP( \
���8���)Om�!��|6��2U^pk�q��� ���^�{g��E��lfSTt�Z�����_��/K��u��9٘���Ŋ!���`2����Yp�ׄ�y�<��G=8�L��7#�����<~�p�!��I��`6���5R�8`I��t�Ϛ�Χ�)2�Tʆ����v�R`��6h�M5Ь��|�H���!:�sMϟ؃�9����������"��+��\��`Q�]_NQ��L64d
	��]��&�HgX������h,il�x3U������x��rBI+	UV�G��.Q��en��l��"<%sQ���/F�x�A� *3ґ0�l�1Z,fCc������+)젎l��Lu�ϓfu�Ӷ!�U���e����t�x>�?��	�����ܧ���8�J�'�W�+h63t
5�\�rD<A��lq?0�3�G�:�{n����ao⌴,t�+�"(���^3ۨW�uxE��"z4����j����ՋMQ�,�����nq���{�@N��QP�����r����G.mEc�[�J��ˡ=t�չ׍;��.��~_?���j�ڸ��~�.#?X[2��n<��g?�t��C��f.�3!Z�8�TI��&�~�4��Q�ܳ�ۙ0�N�����pF!��?Aݫ�h)���UY2��)�s���1��N��Ecy��f�����4ר^�E�$���h��F?���w�U��Y�fy�;����qĢd1�^^��,�E�����{0���n�te���~�nԳ�a���p�n���]�]��76��gI�of���&ͽP�M��8@."�M�ttϓ�/^3M+4�C�:玠x`X�K�E&G�����q�B�d��!!��}ttG\h*�\�b�<H�ϼ����ڗ瞷ۛt�k	f��5�����5����e����%#�i�BR�؍��E���H���!�ɕ������ho��Ӧ�7}��L+����%�Œ@]������ۇ��f���x�T�1���p���x<����\�/p�<��lw��ճ�ɲ$r\6���ȗ��$w����=-�O�?�9����n��f���tл��~���W�gg���ۤ	��&)l>R�tZRKLe*�Ӕn�;������eItp�钬����st!U�)JBQ�}|V�Lv�zT�1�v�i̮A�|e�x��^�l֝�:�?�n��sF���Iӈ1�7.��"mœ�����gn����Z�C��6*�ڇ��}�e�۾������/k������}�I�Ҭ���m��
~D�`�����9�[:�~4no÷[Z=<<`��9><�<:rF#[K���J�0�OWr�d2;�����q;L�}`�~��;��3�|0��$w}�D��%&���i*�n�Q��*z�����L�������HhX'9��a�_K���L����u{����v�F��v�n��!w�k��8]��s�3�����'I.M�SLY,�/�G��5��i�n�m��q�[�7�t a��3\�C�Js��}Ҕ����������ٿd7�o�׳]��s��f��}���.۴��]{���]ϋ�8FX+��Z`d������7az�����Y�������l�K�̩/�g��=��A��$�,۲����{���v�ϗGv�O_�L�1:FC��S�ϟ7������ۗ�˛����ry������[��7/wK���������}���fw�z΋�L�iw�%�:=̄n��M�F-��^��y��̷?����#���J\�l����;�\.g~��R���~����x�[i��|X5�Δ�E�Ywy���a�z�o����W�$�ޯ�{����=v���(��k�޳���~���"�]f��#c����|�ׄ��_���w��%���r9��|7�#N��/ǯ�)g*|0�>�聾�����,W��>(�v;����߿{������NSY:o��ɒ�X��'�֏�������--|IS�@��Z��MF�i��Z;����2{y|��6�F��9�c��!��d7a=O�̎��l�y|�~���@�;�X��|��+d���@��5r���Q�_�v�]r��?@��(�9�|������*-1)hx�����_��0{��$��=��q�� h�b/�P}�,�O9�7��Ŧ`\���w���l39����	��e�]�.$BI�l�7y�����+�81׹3��@�.Ö�L�f���8z�X�N�7�����͠�t�"�]Y�'�O����ˀҹ���Y����|�·���|~B����<����B���83Q!a����χ���kO�~����m/5�=��{����H� ~i�v��&�E���/J�ơ��H���^�����v?��9�z@g�?g��d�{����
��AH����Ұ����d �]�k���l7��8�;��0����pxΛ��Z$>:�gǵZ�����KN~�l����������� ὜��6�At�2�����G��\ȕ��*]M�9R�6󼚯��
�y���V�j5���<O����ρ!q{�x���1�9��+�W��i�:!C���
�� �I��yӜX1�N����)��D�4�C�i��Su:��S{j��T��M��mZ�z��+���?ᬶJjU�U���$V�JTd�	EM�e��y[��k�:�t��:%ZU�յ��E��8�b�f�G��</::ď���H���f����bCdq��d�5��tIO(��n6<��SF�2��D�*��N�F�*|+�F��*��A|@@32��X�������N"�� BM�%H���d���·� *s��<��.��$:9[�Q{�9eT��=U𶌡V�%�R���n��kt��U�T`�T���T�E�u�O���]G������5�ڔn��˔�c6�4�iU�USṴ��iU���մ�>EV��ç�h���k��B� �q��p���N���`u����n:z)3����&ݓF[��+�Z��pA�^Rɶ�=��#�'��b>�>/��L*�r�s	y�RPZ�9�`:�s`�ƔIEт_�[p����[mKHQ�H`�(�eY�V�ʕN�b�~V�J�0✽�iGC^]JG�%d�i��C��Y2�ZR�0�h\���2>
 �Ţ��Zꞃ�ҰΤ86ȣ4���a�D�o4*�i��\�C�ҡ�=WW�_�{����jٴ��`�$�T;0^B��"NEcWܞ��Z�j��㊓�k	t��ξ�Q�CR�W��+ͷb�%%�LtY�j�Y�䠱�.-���Đ΁qlX-K&�@b`D�$��tK�#�kU*�� ��X�9�k�ŏL1:xv��B�C����X��A�x���$�S!���O];R���/C4j9��Ņ�V���֠i��!�OB�1R5ԍ��kz���.�y!�E���:�&О�\	ju��B�
�Y5r���5
��Ny^�С �	)zZ�[���2n�kA2%wM�;��^'У�[$QM�P���u1�H8����uĠOd�J�t(Y����d��	0�s��Ǝk�~��#ژ�OE�[�_�+�G�g��0��/F��JH���mP�#GjU�K�M�7����+ݕ������@��9����drן�
`�#�B�|�&��P���D�~ӽōJoC\��ף�ׂQ�]�T.����&N֦`c��c�8�DsL��ϕц�eAj�8�����Mj��}�m��"�Dc<T��Y��l��l��
���$_�����*�Jl�$�;1y����eJR+Z�IHF%� ���OCBphB�	��M:�R*+!�3�]�f� ����u ^�;�'z5��XN�(�7��aWt��q�
/�V��0t="����Ǹ��} s���8]V�l"�j9x:Y��b.��)�G�JOPV���*AE2�����s��Tm�V����i9މm:9����J�֣.-�8�PH��L��8i������L�wwS�{y��6��q^��6�(j���2��@C�����s�#Ǣ0|L���
�Y'�4���D�`��&3��hp0,L�����=ߥ�:��lɲ��Z��s�n���Z���sz����~JO�Oe���q��W=t�������}��\w��0�� ��`�# t�?Vpk�=,��Mю���\G�'�j>I��=�=�:��H��j�!Ӎ���1�y��>�T�g��vZ�* % ݮ���R�N�nV!v�/��s�mظ�da��ʑ�}�silʁ!v݆h^��IH~�ɭ�V]X"�~s�cK�T��7�'��$:&.���j}����e����� ��] �z�n��`��bn�RE���"]=˂�083�iva�sˠ3^ǬC��"��[�UB�KC��꠯t�b��Dx́O�c@'�/1VaO!����K>��u6%8����w���T���6�!�E⋗�Nc҄�˶��f����$���~ʊ�	��Hٖ��=X슶��Opzg6�����R��lb��o��iQ'�^����<�{�@d���"�.���)�u�5�p.|��Fga�%ԗۜ��zӱ�,;|.�p�N���Z��aw�{f�H�dҎ�    IDAT���S���ό��jσ�����o�1��EX�">M2���+z*}��9�Z2�s$�hwul����9�h����TO��C̞Z��;%�)��ڟ+��z{��`��tnH����#Ke�]Bz����y�떢����q?3�*�"q����矿���D{z�5���������:�Y�ɩvd����m�e�����*�Ā����[�
R��_r��-��z�����-���d�>8�	eǑw�]A�=u���+��)UZ�ǡŤ6��'���B��d���ޔ�>�_ݺ]E䩄��"E6d���K!�2��Q�n�CK5�>�eւ�p�P?t^o*��$�k!cI�����̌K�!��uo�xw���-�y������fd�˰�Jk8s�Q�A(��l�6����|ǋ_��Y�:���M��\��:�b��1�k�֣��*B��K�˞yt�P�;mT�QB7�Nu,E�v��W위�T�bvj�hw+q�l�--~�t�{�l �5,����	/ a��K����}�٬��׌��S0,aJ��)��̥�Յw�'���	)b�����<�t�l��̸������eJ<=1�����:�WX ϵ����s�P܉��s.C~��L�w�t��mr��DMn+�yV�iK�%�Q@�x1�V<�N�nΜG�kQ��"	��?=�b���������>.b�l���l�q�<�XAЛ-jq�.��E��6�L�Dst-['?�=���eGfsi˨3��jj�h%�PT?؉5w�o:SЯ+k)�c1�~Ul��m|��2����x�:0�\��*㾼��M�V S��B�\�4<�.��v��+{�%��d=,gʢwR�@^ක��ɖ���vo�t��\� �NFJ"�f�L�JCil���Vd�����,�Ι�i�4�9w
�]�1��L�v���X"��m��Y�����r� \��k������0=�����zNד���"9����7�t�� ��h(Z&�غB+�����_n��O\�Ge�q����1�'̈�f<]6��B�ORȊ:3����'m�k6�_����Ą�y��}�ra�a����b�����wǇ���ّ;�#�D�{Ŝd�A[= �u/^&j.f�[�]��'ϝ�J�����˻�ݸ��e�o4�*HS�%^l�$zȥ�)x/5v��/�J�Xs��_?�C$��/���l��m�*�cEXp���O�T������x̌;�;Jw�h�Ƿ�o�{9M�Xw��n�Vp-����	�SX�9�[���
b�5���6!=�k�PU��J�$�$�'���P�P/&��1:9�����
�7�6����(��Sn��X�;8���w]&XT���kU�V�F]��-�M�v���b���vzf"YFtAY�W)���T$�n�\�A}�����W���-�;c2�{e��v��u)�Z����G���ڏ���S��	�t�}������8<��gn�J<l�6E�fѵPLج��*i��-�>֎N8�a�%[݇
�%�7Mj��z&C.8�=+��>J}��V+r@$+>/����fS�_v+��6���\w=Z�J��?�Naxѵ����|�!]�ZE��b�w�'*W�s�M@�v�����evN#>	�7FNӅ3j���+����m#��������?�GkR�t:��q�/F"�����t�d��t�d��R�� �s��1��ٚe�	Ň�5$����<s��jw��\oJZ�U_I�U�"�`h�*C1��kq����ﻤr.�/�l��a�95Hݨ���h�o)�����
ĭd���!��b`�I�I@n�d�֋֥*[h1�n��E�C܊�#�G�������f<�7?왾x�Ԡ>O������K������� ��x �8�t=r��B|l�O�ۯo�Z�ې�V�������by��J�[Ɔ#.V����o����%�1�%����JrV�F������Ɇ���x�#0��[iţƽ�^�n�O쮀[W�wM'�+z��Zm��s��>m���Q��w��]�0*]s���i��}O�(B��.��Z��Q�!-m����k7�df��t�RLCQ��|��N�Be������P�X�Џ�n@��������t*�F,�L��@/(8F��UB�~g��D���G�;Ƕ���z�i�nS��,G�R�GJr¡�G����E�@��;Ν�rLc�@U���U�g�x��؊� �Ԫ�Pʆ�'�v���;�9�#��d:+�%S�T�!a�0}1F�Eo�����>,F��|�^|h���ؿ��5C����Wu�0���ŋ��[<�9ϙa����Jm�P�4"�O*�q���hP� dh&��?.�vR�A�c���-F�ƻ�:��G���&??~z~9�{Xo���[o����׵jtP�*��`���3�rP�J]�I�
i,W�5�FQ�Ԭ|MY�>εm4f�|>��IG��Ƈ�VfDw��>3x瞬g�_&�~�$e�9mo�!Fl�4݈�7
�G�VE�M�OU���J��#q��Pq��A���
t:	8RM��l�i�i���o�5?�	��=�]N��w��a�uNTބ����y��7���>������.����םu߯k]�axmb���Q����o_��@�)�	���cV֥�M^Wz��@�M]K��`�y�.8�5�f���9�S��z�Ez�ub�V\�ǝ��VՀB�S�H��h�(\��7�ra �K�3��,)z9/�=.aK��?0�A�T����7����T�
_�cEo�QrЪ�X�;��!#
�plS���E�;��B%_��,�@6Fs�$d���^��ߝ�w43�ڧ�=���Z�>����i����"��Ŭ�m��2q���i�_G�Jr'�'˧67�mޣ �ˊv���q:&8�l4�Aw�a�m��H�-&��l����%e���F�0��I�q)��"�v���i�9��QgD�|nР���P�F�-���O����-���Z�^_�6��WB���6(�-%�n�� �f��Lӑ��;���k���/��|�M��z�}��ƺ/���|o�3�E�kl� ��a^��o�AHb�ꜥ.sg��LZ[Lp¾�e[_`*���4�14�t�Y57�:�5O����p�T�ƨ�Kr.���#aO�mł��T&��Pf8?aU�f��@ ���_ܤ`OD��ZMǋ�	�3��j䀚���/��ː��z�2��m�"����c2�����$4&щ	�s=|zu�<�T�n�{�f�늁^;,������t������Ɗ3S2�)�ה��As&m6r�)�l*Ԇa,ܔ��|��?�x�fFS�{���5wT�$�ɾ�$�ՙ�jz�ժcƩ,�~�z.������Q��
�7�j��)������+�7r�ʶL�u��)��a��m���܀>�c+l� 	`X�c�̯�%t��L�����2�Doh���Ŕ�03�D��z��A��7��g�T/i&�덮�>��_W�>�ZӦ�:||yy������B=�d���	�wEP��M1����$1p��}	�[��d*o$��i�C��=�vb3�T�KW<��P�ɯi�-v�B'-���~@h�#��qVP�&EG;g��P��#�Q��Hi��B�JFk��h�A�cP��N@g����mU�s�C
�������u��1f����������ʓ���&�1ʝ��ͱ|ywz���e��OV�}��t�a�5�ԫ~y~:]޿=��"dCbJ�8��jz�N�M3�d.ɜ*�Tq�Ը� J[P�[��8�D�v��j�%����E�ފ�ʚ���n���^�L�-��H*f���|9k��¡���&n0ǋ���ujqcc�q�*�2���0��@O��~���R��������P�ML�#���H·��i{Ǎ���?���|�tX�ݶֺ��}��t�q`ݞ��g�ˇ��嗯�C�dۓ2r��B��κѬcp���q��) \n&��UG��9f:��(�5�<#笶�[�*�w���}��������bdN�Xj���L�
�c	��0�+���y��ߝ*z�ӻ�`�C�N�+VE8���JOLߑj�y�� `�^����\��ͼv�8��ц�*^N;���#��9FX~��ͅ���N��o�>�Zb}�_W���'A�t���J�~=��K=9M��L��<:���Uoә��Y����ð�U���V�[�W\ضq_�#)���9���ll�z��?�բ8/4���S�����)J��$�:�lc�x��К���6Ѵ���NÊv�d7U��&��V�+_���20�|m��L�jV�ʙEK6�t89��v�D�Û��~��`�n6��w����"t��0!.�z�������?�>��<R,����ݜ!�&
W�p�8E�L�_�Y�9Y�
�w�6��V�b�୲m��U4��q��4�{<#�QD{'��{0'�nc3��{W�0Ί����?JՊD=�V�����a�ǡ�ڮ[��8�uN<;�3�QL��0}����-t�ք���+�L��8O~uL�QgX�a���6Z��V��=kw�}~y8}�pX*0؞���~]�F_{6Ӹi��Q¹�����f՟�Mq#��T��Ɗ����lP����1O�r<m�Ȋ�#1��oB��"�m�a�\%�l	$F�=1��3�V*�iWE/�1�� G;A�4���ca����y��9a��R�4�Z�c�; ���&������I�S#;��G�8p�� 0wwd�o�o�sJt,�u4����,~�1�m1�����p*��E�|����pyx����{N���~]��:*�
�7�_?��r��I�ά�y.PO�����	���G�j�թn�7�\����}�9��`B��Hi�YlPP��Z9F+�c3-�0, �ZU8���4�dhg�چ�[?�aM�ѱ�(�7�ӱ��S��2z������y�f�U=���Y=�`��=�j�n�D�7U��1`'��_X�u ��w�1�.U�E�NH89����ռ�޾P���������.�ٯ�]�=ֺ�Ļ�9������������OU����7��k��lJ�%U%6�c}kD�x�58�J��X4�c��)%�:�K' ��Ҳv���Q�FoJ�'A�Z&=jn�8O�Zjn�a��cP��8VTrMey�?{W��*����^�P��,��4�D�Ĳ4$[�H�M��I�鬢{)O�?�}�!��?�U�/�����Ƕ��PpQhx|E����� �����7��N�r�Ft��6Bۖ�5Z�1�����5�M���˥(\	�s�T��b�M���-L�IDKY�L<�����^��G�X�z"�F�=���]=��:U-��U��i7�ů��*�6(���r�̵@W<!�{�q;jp� Ɔ�A_� ���D�PPt8�('<]q�9�o��F�󡖕��8���T8ђ�7����8}x��>}���XT�9}?��!:hP؃��m��@��9E=�i���9(������?����V��و�H�J�B%�����HiU��%����-�r�B�}4�V�65���{W�����ZS��ؼ���+m���&ZUfb��{��7:��/�������>i��<��'�x��i�
ρ'!�|���^����W��f��.E��I$^xEPI� ڠpڠM`�o�޶IK� �d*8��.�$)�S�J���2$B Iӝv>^�D�������C\�Yg�)#��>�����3��Ԉ�z���n�5��ˍ}B�ǽ��{����0��x�9�ޞ�n�j���ڝ?���?����n��so�^i��x��������w\���v|v���iw �N'>���x�7��
�̛L��c��vx�n�������t�Il��؝�7�ӡ�fs<�d�H��#6�x ��ԑ��	>����p#?�}�H^�	;�a�����~�QL�XH �,��� ����n��<���͏w�G�`��~_�,T��+����3xBB7�7z�2��l��u�//��"�/��~�7��lY�/��Y�zI���u^����Ҥe�T�p�{��2��r����a����eZ¼oh��9��ͼj�y�xJbT%��eS6M��y熮?ĕ��z�'��)̟Rz�M���:O�u:_W0VUU"{5��E&ҲN%0�R�F��DĬ�����uY?U@�Ó��Ҵj��F~��eo^�� �&����7os_ί���^���M�I8�)آ����\o�����%!'\rV�8�bXb�1�3:���`��Y��b�ӂN�\t���n��t�<�v~���� D�>Ѻٳx!�.�D�}"F�lH����̛3��G8�t�c���$�.^�2�Wޱ������	���Wʳ�Н/���ɭ!-�3�|�w��}�E�C���gʋNU�n�#՝��/��e��E��L�n�Z.�B2@���|��"R![�77!9��G�8M��J�����[%�a�E�0 ���@>_�;Sd�M˂y�CǷܬc�1����t~���-�(��Q��?�}����S|p<��T���|xT\�v'�;|����+�9��Q��i����W��7�(T���Bo.��.�g?ƞ=��q�g���>o�}�4%,���ْ���;�v��)Y�|0>)y���?e�V�H�o�OU�[IHAs\V� �p#���8(U�yS���0P���K�稀D���p�U����6��G
e��R�|_^�ݯ�k�*�1����Ev?q�v�)�US���r�n����W/s)"���~�,�y�� 2���wY�_.T�)�/u��{�z>˛�K~�������lȿ/�de�;v���Q�֭���4��(��P�u)��7�c��QF���� �^H��(�C펂wT�E�w�Ep�~�) �=����۱��Ķ9�D��=�W��y�2�Zu�U���ō��n:.�,�2����,��r�w����gT�q��A�У����÷�;��ђs��~9�x^��"<>�Ͻ|�2e�i�k{�n{�����ζz�����:��F`��=h�6�$��N�9;��'��$)��M��p8I��8nEE^��v|s��s罂ċ��a��D^R���	�H�؊��L�ɼ�$Nĩ�" xQp�S�98N�%Q?C9�۰ES�EA���0@�l�`0h}�ִX\���>��f�;Z�b��)z2�XǍw�u��4��Q&�vV��6���̐�)5�����y�~��� �H��I��\� �����Y�a���C{:�i8Z������Z���r��2G\gJݓ���!�D-5��
�C���`�]w�WMTh�D�kje��zT��>P����g��*�i}n�����XY#�:�<��,�5ؠA���u�C����c�Hc:�p0��B{������j;FQ�b:J��$
Ѱ8h#�9��1�ߔ��T��?6�,iy�Ͻ�����^�Y$'e���h����45u�@=CK+�K��A.K�d�>��E�M������<!�.����K���\f��L*ڃ��a��Ͳ�adCF�H >S��JpU
�j�!�H���U����u��0���X��Z���%�k9yJW<��PJiFJ��w�:��F��2)`0
l4�;����@obX�va���>_i.�'�I�;;ۣ��R��˪s&�C�nIv����m��椑=�t�p��ˬ���Z�Tl����Xj���x�A�@+@`�d}���^}�����������sm4{���e� aT/f�nM���q,���O��sԃ�\�5z�ʶ�
y�N� �ԕt�'��V~�)�
_ �y��`u����C�D?J=ʐ�IW4�Xpmd�f�ϑ1����Ъ*�%����(���Í�I� ���_��KpR+�a�U�#ao��#a��q�j0���6�N�a������a� ᔽ��r��Qw��4ZeTT��'�iT�����a�nrH)�v��a(��jA��x}�k����pϾ{�_�s�:�'�)�]�Z
�/]������>���)#M��D�ժ����q*��
�~hVzy
d���[�"3O�bW���.�!��r
g��\<kC�x��ob����{��ZTn�QK䜱�V60Xf#8~�X�r��ӏ�t�O��2�n�f�>�-���])�+X̎��*��� 7M�T\'X�R��z~.��g���7J�
���n�����5*��mL���7�ɕ��נ3��ˑz�zs�/�_0�T	����+M"�z�К���X�:C��F�����cu5dh��9$�R6���i�1aR�$˿y�gq�P�Gdf1A����d��y.��VOM.�W��r���"���� ���b#�\6q/���s�h~�_�Ag��('���ߍ{p� ���}uA�j�pyW�[:�T�>t����q�bg��X������ 4$(��p��������?�TQW�ل7�\B���_0!\a��ҸR�=�ߋ�9|�ճ��sŭ�F�F5�o���OG|��|��O������Q{}wkuG�P����(�ٴ�!ڲ,��Z.�+z��WP�Y�r��Q��( ɲ�u	C;����P�{ܺ.��lz��m��啕w��Ŷ:�AC���ڍ���0�_�����c���	x��v�t��e1����X�(��A�Un��DQ��b`�j�Vq쉺��������_Ds�z���i\Ȭe�;�Z6�	Bw|���k��v_B�`F|����=�ȣO�;wN�#�B�kQ�<d���Ӓ�$&��)����#���v��w���s��j�z��9�_!C�&4���p^6���yg0���[���f��I4e���4�����;(�ձDد^���}����;H���������I���i\c�:��Μ˴Q��$u%H{����>X��B����n쐈�_C8`���Z����)�C�C��8�6����;��yC��5φΗ��b����<H���z9q��h�ܩE*1�U��X�0��6cnhW��
1[����U-����HCf�ѱ`�?ߤ[�9}9����n'��W|}�P_*���tj+���bab!���p���I�?����Mal��f"�s;�!�H�+5�1�F�z�bx�����	֯�dvQˤ�RA����+��=e�3�I�,+4�oH��oT-��/�/��J�ݒ���G3�����p�o�٦�}��K(���G��&�n�|V����ͪ�w~�ቌ�,U��*����vG�������6ޢن.�̱�[�5ueX�P�%�ts�"y�xt:PdI�$I�GHJ��B��,�c��+�Ɵ�����5"�3�*���j,��Vc����'-�o1;3
�>ؼ�C�镍^Lť�X�G��S��c/:{e�J�q�v�6`thbq����HUH�oi��:�|��4�6wۋE�*Y^���]d��-Ŏg*v�Ga+lYo��Cm�����=��"�6'S�߭knJ&�5�sԑ��tϽ&Sw�fh�f	�N߷Z}Lg�fo�YS�%��}^���_��T�e��q�Np�n��e8���!ٶ����7̓F�>�,W)�Q-��[��P� �hYP��:��QS��,�������~�2Rt,���s�h�ݶ�_;|�-̖��yf��q��ux�ۮ���i�_u����nL%��?��
r�]_H|������q��:�}�X�|?��mC�.=�+j�2q,�­:z���cC�L����J#��r�������&5^�R�iK����*��<&���f��S�QGa~����7�Ր�=�:F���!���4��P,��Ou��p���_��1d1vj�h'�2��|�
{�E��S�V$�Μ�kv�4!��_���g�)�#�V,�5��֔7N���Q/v<i���?�ʄf�_1n��N�m��o�T�gk�F�ⶢ��g��1����pӆcɹ�^,g�l���+��ۤʵF'��}ݚ%1����p���NЃV�Ƣm�����{k��n�q�5q�k�)��Y\��o-���-:�"�ٯ/���{b���\3��w	��ڮ�晪h��;��ʖ]p3�M�y1j<���BMcԪ_&^���Po�"B=���I ��6g��ak����n�Yf�<iݪ�5��;O+�9�(IX���e�-��wR�{�`t�:�>�J�g��L}�|�W�|��VM���T���D���M��j��i��z�������ûOT1W��*�ZmД�S<c�����a�P����v�A�u�����`����r�T��V�9�l�~�"%�o'����Fl_ �nuڣD���6�'��Ͼ��o�Y7�t��f�D/���SuAc���}Y���GX��U�{l���Z�j
�:[p�X�1��YB#=)���
TX�	؛a%�����N�p:��z�8�guOSLSz=�g�0:7u�WF��n�i�q�L���9���]d�_���b�:����J&: 
Z��o��(ga�����{�W�k-[��I!�S���m�/W����[XD��(��.Ѽ��d?�b���f�xn��~F� թx��L��M����2�){�6����yhoD�==h�b�-=��^o�(�χՙ�a��w4��`��痭�7�UU�fKq�K�����]�Σs�%0ҦP 0�Ҩ)urѻE����<�Jk�}}�꼴�+*�j�"K�*���毱ӭ�#�F��xL)�I�4���"ߌף)s��J���v�XX�fxw�����2N 
F�[ʹW��kC��{�V��l�'>EP����3&���ш�"zR�7H��ib`_g�ǿGS�a=�䗤�ܛa�}�Z�'i1ȃ,�3ߏ���F������P3�����\}H~b�jm��`�.���c~�_	�(���[ۀV/���c�Μ�E���3ޙ�ٵM_��:��R8	��a/U�F�o�ߩ�^�c|jg�<�f�Y_�P�<E�ܶ͜l��?��/e�%>��N��~�i�_�����Z�~o�`��X�v�a�Bv��T����	�1ftɧY�\~�C��B��a8Ãa��v���������g�M{o��ٺ-��|��A�sog�l^��E���� Ғ�}R��w�bnҡ�'��O'.��H��B"f���5H$qen�F��N�v��5��jD;+>K�Pb�����s��_�*�Ȗ������	1h�#CĒ��H���U��(�w��{�|��0��]�C��]���ދ��yK�%�������Z*��1z��%�7P��
�7N�%E��E�[����w�$	�[Ǆ�����#��P_�NdyEܟG<u}h+��q^L��GW��6�pB��"Y�pk�D�R҉(nk�(�N$����Ou�Yo�^�^��x�D����SD��dd%_X=�W���0��啫��v���gҵG���Y��c炖���a+GĖA��e�+���$ح~�RT��q���G��N]�m��6d��aNb	�[X���p��j������tKYٗU���iQk����"����8��+�R��V�����p�O�t��b��@)�bD\�ӏY^s���DBtf?.��K��#��m�O��%��d�V�@ 示<x���"��m�:���,Fy�N���3 Y���1����tf���lk[�z�BN)|���v���T��GqGaJ�Am~']W5����v_|�xyyhꗀ,h��do�S�R���B����ab��+^\�?n��WS�aT��s��}�lq������Z}\��h��d:2�Z0A�̏%: ���.��D,�n9��6A�ΰ����|(�ob	?��=���ɦ����vp[�?Wgxt�պ0'1�������)�brF��v�U�ߞ:�\��J���(����������_7_���6����b!6�*8;�-����>����Q1�\���]I�o�*F���y����~W�W��pA�]W��Sa���0"5�=d���R��F�*A�Q��Wn��q��)r��b����*n�m�M��{��V1�8ٌ��n]���+�LC��>���	��i^%(�[m��װ���X1l�+tIx�B�I�(l������C_L֏gؚ��͊%��I�Y^����}�M$�Σ_l5n�?�΄���#M�)�c3ّ�	���G.�bf�U�뱬��xvEC)6��v!wW�djb��r�[����Jօ��*E��~]���tH5���d�ރ�������h@`���u�Ɯ��?&S������Y�|�t}��Sۢ:z��(w�Sn!q���\*^��m/�^��U?+���x�\%�[Í��d�T.t�&+�@SL�!���G��s�~҂�d���4��!�	&�(�8>;�HI����kb��-�c�[�&�Ye��}��a�3ɴ�e��̓4�aA�a��1��Y�,o�d�l�q�_�d7P�&pHY��L��dS��%�V��pq;��K��PA� 3v�F���X�.7֜�tF���Rr.M;Q�q�b��xN,�@IP�5ˠ�F����^�����A��(�ț�2/�<�)u :@���pߣ߉�G��]�.��&���T"f������Zc�'����4dZ��+�2�,���,������}h��j
����4Q�ps�*��.��s��ɞ� m�{�f�Γ���1�:�&т\�?����(h%���*���ZLG�&�>/6�Y3A���~�
�n3��`Ev�F��NZ�@2ƾ~����W?O̬��������Y�^n?!������7%12^���3��-a L(���O��^Gc�_וB u�A��e����ܭ���뼼��`rPT���1;I��a;U�@���0�-E�����~�S޸��2�xs��+��0k^cUA�z�i�<CPs�N����8�1.v�~��@�	�ۨ%�EpM
�B3��W	����n�A^�t!�Y�"���!��ҕ���:���DZ�Gۂ�ɽ4���x]��G��}��g��$��Z�Z�O^�Ը��l*���lW�'E�Ҟ	Y�bv��~�9� ��)���ߝ|�����mK���>&D���<��P��Cۥ�D<�(,N{6��R��`Ma���g9�W����]Fr�Ȁ���"6�����4���9s	$k�&���a0+�U����^�=��Z?�f�F�Z���"���|���ÑX�g	}���5s�?'�C����l�[gJ-XF*�#���痠�/��g̙k�~��7���R�"��Vk�jDܡ渷��U���}��}��0,�SR��?=�"���w���,mr�y�b̂n���2��ϫH@�o՛�������%�%���%��[�s���؄�����B� D�Y���?�*v�����D[f���뇛��f��L��аF���j�G��'�ESKY�#}�_5HO�ڸ��VI^U�83Q���%�Z��i|Xu�g�����׫���ٰ���QI�Z����G���\����r�)iv{9�R�5���2�J�SN����h!����@��r�0B�ĺ��g���8���f�9�\`nנ��a������z^<������V�F8��FA�QbsC������冉ĺ���ey�l�h�������|�e�zqp��=� �[k�(ՃDCD�N��i�>1oks����D�,�~'�	�;ޝ#_V��6����w
��`�8z��c���+�T9eU����y����<�=R+����b{q9�P�N!�RL%jaR@��)b����+1ס˰9��^�B��h�[���,��"���O)��p���3���x�)�J��<������g�?��X��O������z�e�a*���f�,���AD*lb�Mʫ�uL��؃��s��;�5���ߤ-n7��b`7���zA�q��G��r�������J���c��W@f~T�w��M��3����H*{�����D:v�~���+A�c�P�g@�fL{K�p	��<�z��ѡ����Q+�����qǣ-��@����i��8�\ ��2�<���`b����+`!Jp-r'�o��ϊ]n5�X���7����]@He�K���\DN"�ݳ���V�*%�l��99��q�0��/&ғܽ��� Q�'Rp�x�d�`������m	�%G�^	��:f�)Y��3���,���r���<�4�'��(��F�UG8-@p��`����\�4e�F�`�c0.*/In�~�DM��6������S���E�=�z����Y�+N�Bj�"K$f6_j���P@{�j�h}�T)��eI�1��ώ�������"L�t�[��?�-p��+]<}M�1��� rIR7���y�yF�C�^뵇�ߵ�z��m�	ȹp�\�~ ����Ɋ#/ض�_9�bǔ|^3K��=Ҵ-8_ۂ�qt$֩&Gmu��������V߲�Ȼ��@�������'U6;Ы��6�)]������NqA��qe�������pz� � |@f��=RvH��70��"��a��"cM��c(���0��J�>Q����zA!k|I>	$�}լ�y���n�*ge�hy���J#ul��h�o�S瀘�!�=e<�������l��X�_UT�c--`t����=A�1�X����ް�,룏4�)����w���zΖ?��8(%�t'M���c�0��W�� S%�>�kH�6�ˎ.����;E�2u�M��DZ�<��!\w��{=7M�I	��;��H��{(�]ﺘs�U�}%H�}���Q��uV�9��?8ָM��	n�ڱ��=P(4���W���p/Fܺ��8�t�>8�DW��?R�`�XexY�a>����A�g9���ߺ#�wu��u�|>�ύdH���M���-�K*��\�|I�L�ƚ�0�����%ʪ��������+y?�z��;G� e���3�P2�2���H
a@>l�0�ZΉ޺L�Bn�M�p�\o�\�3�GQ��'���nD���N����k�:�5=�Z�XW~#�'R�kL����)���
��1pX������
���9�6_�
9>�!d�Xy�MR���)�梧ԧ�D��m�������s�����A̻�5vB��z�k
��c�Z�0h�@<=�䊦�'�����+b�P�b�;j�{�ZUJ��6_����ZPNn�K��=������.t�o���*���8�1��//�Bd�E��U�L���2�z�z�fxy3���L����0��Oqђ�		�H	X�k���p�Y�=�O�<3��}V~K�Ûl3��q��enQVCr�o�ز��˭NeNE���0�̃@d��R�>�k.�>̐��v��W�3`�:6��)���0�ݯ��\K���K�4M����A�����9�Fd/�*���uã��C�={�|��Ґ�%lEg���3�(x=(�~t��[����ߦ�m*Y�G�(���

�]q���mǻm�("AZCQB~|�rcnuN}=��%̠�|D��'�X���k>�'�/�	b�}u���*�Q+>J�0g�ڨU��{؆��Z���wp�n=*�_���ߖZn��`KJ��Y�����N(�L�
�����c��ϘG$-�	������7f�0�!;����a�s-&Jcwą?�ﴄj�p;kj��U�}uEpԚB�{������΂����F	�	��N�?S������k�f̷鋓X	��_���5�6��(���R<���Mrfc�J�izO�t�栩߁6@�W	W�6̿�J��g#��0[���]ȍ��m-�����G,�����/22��s>ԗ�+jY�%�u�D��i�·�����l��x�Cf�������5`ɶ� �yW]t"��v"ei���u�����Bx�ƹ�zp�"��^O?��R��w���89 �i�d[H_�,����h����E���L��`�佹���}@�~���)%���C	o:��W��.z����{����kn�*�?١��=�����0#Uh�Oo��oʌp�5��>mR�j����z��(�ק�\׆K���k�8'C�!˽�z/3Aw~^]���D��?������-u�P���] �pǲ��&��(�LY;o!r��*��4��LM���'h��{�m��������O�
���Y��Eb�[��8�Y���i���$Qxk���4iH�Vem���!���־��=?�]V�}պ��L��-M\�5b��YGp��\�fX/)%Z�%](�sǊ��'M�9|�xpڨ~��ӛ�4����
�Œ-�dsƮSwm�e��E����/�Oaē�;z�v����)F�SZ�Ȓ�48e���=���I���,��J�Oe�#
"yθ��¤�|VZ�!����uD*�^��
q3WU���D�����a;4���e�"ƏAZ#O�<[��J>H���CZv�LWU"��X�O�7�s���2�o����P�鸺��q!.�wYv����˒V�|�:ߵ�Ȕ��[d
b�b�驹��2k�T\P,�xuh������+ү/]���P]���PLv�d�GOlWhy�����Ҫ��U�t���R��K�d�w	"2�H�ⶦ��ɩw/����8T�e����8[�0B� C/r�����}����p�kŅ<1[�#�ً���wO>��=!q��iY|�uT8����[��e��Yg:��^�3��1_��xXt�s���pyt<��K��>�v��\��ME=d|����ʽhl�IA`�̻��� ��DC5��S9��c�����\�Ph��\�4;dD�:Yآ�-~)S�mv<9ߏ�-k2�����$�<�� ?-�'-�'�k�a�H�L�n`{�!X��6�2)���z���HϘ�>�C��9'ě�3yɍ&�u�L�ԬW�6�����tk�.d���q�hϕ�>��CX��f`=�Ä�?��Η�� ��}���Z��'zG��+�{��trh.�m���2j�O�T9}||���{�i��m���nA�W�#M?I��U&x�� ���ccB�b�G��\x$m�I�MXs�v��R����O�N����n�VX��Gd�n �0r;9@7:e��M�&W�o�0��`�b���̘�I���t�wPoS<��`�`��%�?67qp����}J햚;>?'�puy�,U�;ʩ��u7��<����v�4$t5B��{��<���}��o	KkT���7��)���V�"�7��7���z0bK� ��������!�k�aN�lx}�)V���eI\����Y굚�b9�\ZVE�u�vO��Sm+������339�L�{#��a�%���ފ�Q�������W����N�p�y�2R8ڧ����&.����5�g���N0�_�Fp8pjQ^6c�(�!�w�X{�h��|��a֜�2+$|��:����>ą|^�.��x��|"�$���T;*�wC^���f�v]��"�~��ݑR�վ�=+�9.碕=x����x�|vv�GS-�/7?����MY'�X�>����G�dln>K��|�A�.����Un��q5:���R���\�ޟ$?�&�C6��J9,����O��u��K���'��s�4��f]�P��M)�U�n��57���:&�rUq��r�K���u�ꖓ����lo���kE�jsyV��6��S;���8�|k���٤wQ���1v�8-w1����Q�����=CP�L�%��/�J�c���W�=�*]=(�Y�,ʥ�Rܩ���xd#�~C�V[����t��C�4^�sg:D!���Fq)��a+�|S��z��0��NG��T�6��u,��!�c_�]5��MH	A�����U2��մ��u���a7f�ܰ�iNX+�uP���4�x���?�Tk��.~9�j)=z���M�����.�j��
�Ǻ��3���_-n�dR��d�"���7CTԴ0|r/��-NI�o� �ʏI�'>��:��&��+���S	�Z&|�q�/b.����\�f��-W�)���+%�XZ;��"�w2ѓli��xjԑ��9�0�g���0q��MLpc)�c��%x�ŮxF��]`�1�,�xL�UhD�ᔚ���l�G��+[��}
��gu��
g�P�ϩ�����Z���p�d�P�廜�o:V�R����.�27I���&��ȷk8�뙷T�D�D��_�ǏK�_H\ۈ<�a������R3��H�u�z�����	�e.7�h�J���m�ƴm̬�;O��/H0uX?|�C��&���l�%TSI��B͝,�n-�/�R�C��/W�X��i;$�RQԚ<�]�7L,�W����1�s���1�H�忑˷��q�$��!��&XIV�W���ij��|`;�Yd��ȡ�:%+����N�(�Ol��Ү�=�u��srd2<v�㺓Y%��2��'R���������gO��b����(�b�N0�RYY��D1Mt��[�:�E���-�\���VT%�ra"��b��$���\v��!�*L�³d
���B@������\ɀ� �_ʦR�Y�~Z�;D�Iׁ祥�r���v��"Q�G[�8~�����d�VQ��e���ET��BdޓƷ@k6���g~׌�Y^��F��AI���̨i*��;B�йD%�cO���h]3i��$A����NM���F�������>8i���	0�3M,���p�i8jHd�_A[���DS�=�]B(GU��t�_Y�t�#˺]�!Υ:;+Q�,�JkM�z�-���.�i��}�gHe�h.e*�c�s��l!	�9RGj"�>w��Os��.Z�A���'$�%��~̦��G$����M��@dl�:�Z�&wP��{x��3�O�� %.��\��F�.���>����>�À^�?��Jw.����
V�����Ij�)za!����h���0�j���5��^'ٕ���Vh�S����=�����������K:x��C�%��^�-Byħ8v��{`Zɗ����)a{�U��˔f����^53����،kX,&͚��v�Nl�(Q�+dEM� �s���U<_@��NO�1=�]�}�y���Jn�Ε`S�� �z����CK̈́Ur,��ZE�lgn([)��-����bCv�`�?�I���EED��o�J~�*�����'<o��	�c~�)�vKII��K=>�o�s������l�@��Я������L���B��=�vY�9�vȣӛ�ᬶ��UdNU���.����t(�9Z�k��a�%.��秨��( k!+���j���_!`J�����*v�A!�ef�3����;�����lݞ�6�����v���nC�})����EV�VÃ���#��'{^������]�<�J�������fBG���(hɎEV��_~�n��|D�W��/dɵ��d8ϧ3a����2�o��03�۔Hng�j����ț�k.HT�Z��fxn�!�[����	��k��D�q��ߑ� b��o	oR�FM����z�G��+�Z���
&�u�VT'b�A`T�u6o̧�.�5m���\��[d=�lH�8�lu}9}-��k�M�+a�Q
'X��|�?5�=�#o���>�wX�E�����C��:�{1�� �RgJ��U��"ZZ�cl�5�J�:1�j�5��Ҩ�:��{ ��<��>��L/~Y�����
k{�/�#�UI����<��v#�2B�fD��꾡b��fBYa�'.��{�A$�BӚn`�9�.�� �^���/k��:�=
�����P�CR4I�_g����Ա��C��1
? �mVW=��[��T�ѐ%��#�I�s������A�+��|A1�������z(%Fq=E�	�쿸o��㡯�GS\���,�.0C������ҥ��7�.}(K��SB��E���j5�`�M@[V��c�DC�$iU��#0 ���]
�$=��z���x3L��`x�C�a�<e�0�}rY0	N�Z��Z$����T����>8����,����$zM��|��/�Y��O|��s�H��8��#�����?.ĺ��؜�B=�;gԲ���j�fY���#��Idβ3�25E��H�Pr�k��Zh0�Qt/ <_ 9��WM�R+j��O��iY� �d����;}µ�������)������Jɉ�ïu���<z[~�aO�k���M����_�(P�}��׹+�8�8�yD��v;��=хƂ�Ӛ��گSS2^F{�3��"�W+=T�C{E6x��K�ػ��z`�bG�]U��G���1t)>�F�	��(0q��ז���e��m�L?X=��Ц�a�(�DB�Ю���\tBjL���R3��3f �}���5�!�A���b�]K�����i�6Bx�|v^��.���w��8��������{
���,hXq
	�7� ��8��;��@���O��{!��R2k>,�5�;?���L�Km.���ʞEN,ˮU�t��֜�^,gSvdA��ً�nb>5Ό�\i�;<l��Z�.6�o�6�9��fե��^���m����7��scv��ӹ>��#]2��ب>Í~8X�������7s8���A�'��9��G�򹌿���?�^-��ck�p�i�89dOb.�W�\M5t%�@W�q����K�P[:��˟���H��[��L��ghm��%�,�)̞4��?�W�$����"[���]X�B��������٬�G���K� �K)p�(��Gn8)$XbU�&���	���a;��+.�}d�V蓂�k.�r�wMuK��kwGaC)���w�%O�Ic��ݦx1h��?	���$#Y&D��bL�2ق7����c�h�����y���l�\}��ക���4���F�\yQ���0�H`#�O���؃&7H���S�9��w�?���d��B�\��z���!��7��b�}7��Mo���>��ko�8=�5�ᠠ}��^���F�|)+�~����)W�I��kK�{T8�"S�2'~�֖�R��e�:����>�i7wC��|;�}0s7ǩD�%rYt��ܣnܧDi~R0d��M��V�0y*�s��𗌦0^p�LWAӅE�»�dF�z�}fA����9��zisސ��o�y�H��������3��l�*����X�I��gA�l�A�4ﵧ�0~�f���[�K�p>2��� �k�v�-�����g���d��x��1l�l	�fm<��k���a�Ɗ ��'�h5�	�	�AJ���}0��0-��!b�������F�&�rl���𯋻T@+�ڂ捩�=���z�e>�J/�ȷ\��c�P˝b*]8�cG�d��ðh#�� z/3%X�|ՇӷN=�'�(��[!� �\ML?h��.{�}�3��/p ���aH�,ڝ�ll߭T�Z��wcL�]M.w�N�%=#�X��6�=��9�X�S6�k���,�%�h)��i|�R�ST h��lQ_*����Y�҄���� �����YtP��{R����r�l�vF~��6���\�i�j��/yU��̹���"-����4�䎹M�O$F9sj��d�<M���dվ^f^y�v��5����/���ÌP�IQ�$�NF���T�5�Ә�dk�I����Xڇ*�U.ݛL8�q~��<b��sJIkz4D\؍i"���IZ��m��;�A_�QkI8s8��9}`p$�Lb�q�oBJm6i�04.%/8*g�ʅ[��Ԑ;�#�"�SSH����3E��N� 2�5�-_�Ud"�Y�a�ȼ���MuŐQ*b�20�CoȳT	�BF�� �7����~���Z�l��g&ҿ&�������_�V��毃.U������Z����<Ъ�����P��&HN:hDe`$��1��:"L
�V��M�9x�}{t[����"k:H&��d�W���0���Dv��DJݗ��ʝ���!}�ڞ3U��Ĵvu�\�~V�&e�S~Q����#�j+�Z�r��� ����A2f�Ez&���CК;T� ��\�lb��E���
��P�%)�8��-C�&��l:�ޣ�<-��u�����J��x�tW�����	D;�a~>x5";��,�S�����a��F[Z���b�ek�J2�8�(c��e�gy>��@TrbASM۲Y��i�x�F�t�c�����V��v�Y�ހq���>�:�˰��g޲_AI̻�.N3C?��͆�nz��j<k�R$���+6�\�1���\gOa�}��	{�F��6��%a�R��Y�����o��?��m���d�q��o�����u�*�gÐTJ�z}���Y��Q~�d��_(;���m0��bN�瞔�U�����@��}�f|���Kǐ��0�=�+D��=�f���%���UǙ�̅��Z�_���qDljN' ��OrG~�b{�_Եzt�;v�Ϭ�0$:����<
���V�r��j���J��0�A��]C�&���N����-�	{�^�iq�c��|RH�� l�{�V����~9q�튗u����j [�j�u�ӂ��-���^�Wo�ٕ�l_��eO}��J�2��+r���~�\���J*f�������t�r��c����(c���G��%c��-�9KnH�U%���؛C�� v_p�:�P�4��bu०pK��G�����c]�:�:�!��&9#�����7E�_�L��z9˿9�4�"�*�ά������҅"�?=G��<��Q=���`̀PC�eF�����l$˜��b;�U�6�L��i�a���X�9��BߞD�r�����_�&},�5i���IOi��d_0n�,b#]g9�5X	������I���S)��po��2���[���c��0�
���I�K��>(mr)�oȺI/��0W>9Pt��k�a*�/����!�Ba��f��]M3D��
1�P�;o� $ш�W{��>"~Ҳ�7Rb���}{�T�����f:�� �[��ͫ����������A���_~�P3�p�[�JJ�̓��#���}7��iH�P�~�-�^�$�!\����dUm�C쐘�9X�������L8Ħȱ$�AH<�W�%�n���'���`����~�7�����)���[��z	*�`_l��1\'�����~�/�PV�eX�bc:}�ed�.����@�1�����\��W�uLz���!�[�o��/�_�EMte��"���X�LK,N�/j��g֐ٰ�z��qѣm5Sܢ��D��e��D���р�ڽ~_嬋�	�FIYZٹ�~<��@) ؃�����/,�Uz���n�,#�&��&+�`EPDb܅#�5�z���k�QGې��T�Pҗ?r-�1k������+�����y�7:�[?8/D��� y̲�XE�tE����n�y����hN2�H��O9cz5�l�}�:s�����dv���[7���${�L�A�������Ʌ	�
_������?�b�G��V��+�/�$S%m%����-%R{�ԇ4�;b���gR� ��η9�9�}ѯN���F��U3k�*})�t�:���q/)8���J7å~�x>�/1��w��*��y ��Ly��@ =�6����/`�}sύ��P�\���)yc�;D�BL/�����������q��q>�Wy�ys<�����z�]�+(��!�6�#ʶ<�,���OB�a�b7����}T�sȖ��^'{�D�f� y~D=�C.��y �h������|ix`P"I ��ŭ�s��g���C�v������r��)��5[5�yx)�n!��.�=�h�L����;�MJ+a��j�-�ζ�k��+^��}��g��j}�ˤ�v
��ob�_f#j�G�<��A)�>��tNXXELҒhv�fkd8Y����cdSZSh�����J�~���L27�2/3�����z�|�,pX�?YƔٰN�+�����$�|����s��&LB:9�w!~��N���fK����5��VU�	,��IK�A���~jGW���%h_&o�F�$0-��StT�kZ����A�xPx�\�{s<B�.O�I�L��P͹�g&F����X5�w��[6 ���������'"[Фem0'�~x	���0�̖o����e��E��gI�@Wm�¹�"�a8����3οfGkI���!m�'e�ˠ?��+ԑ#_���pK�/���ѫÚ|�x����5���%SP�tw�hi��N�QR���k�����h���s�k��{��?�'����/�J�Q?�#I����	eS�=4p��m����������	_�,�(�v�9t qS� ����Ѽr
7i����2Ɏ
���-^_K>p�A�nC*�x~����$����8�->�\�e�c�UI5:�N�)���z�q̋��Ţ��2���L�$�wdh|�[/Ut�#ѿ�%�E��KJ�6����O�q��a�z���l��P@���0��6!��EaU����<jKҫfƒ���_�)L�75ƽ�
O��C��pӨ�]��Q2ـ�,��r��f�:a˖�s��$wt0�N2��B䠈�~33R�̷�酇�L�6�Z�q�"��s���Cx΢���3g�y������)�*7.���0@�]�ί ag�������v>�#S�SU�=�qf�m�I6+n8��Y��6�2�K�z
9�$�,�q4�R��m�J=˻�ě�+����W�����c(��W5�m���=��L���[��{f<�ѭ|��5�9wF��j����ħ�R�UA{4��2�n�����exg5t�y=�8�N�Qt�N�7W�K��<�`X�V�V���_͜�\8(�����Y�ԟ�L�;.���Yv]f��0����j�2�G�-���7�-�1�$	���rGJ���h���݃>в_K>�v�Ș�6L$] v0s@s�iqd��yaֳgx��tW��)���9�^Y�O\I�
�.A����)K��(���)��ju�Pϣ��R�L\ҜS�h��%|0S��2ì�㮌Þ�?3pݲ��j�V�kҴ�k���Z��k�w�[&�2 ���\��|������BoVf���������BP�Ͽ��J��F�0�q��(�h�RwE-��� P� ����� E!�k��'�s�a��`�}[c����h4�D � Z�G��%3��uc�%�����G��:��n^�7�M��5�p�����;����ެ�X��z�S��7���t״�jG���V�d[��g��x��!�t�Y��s�|˄�R�UY[�����-�3H8����v�)/�1�nx0�[�Gh���7����[���Y���禷Y��eu��|R�� >Ky~>���0��}Rf�H��m��aI/���?>[3 LT��+9C���F��YQ��9}�p���T����6�Bx*���)������<�$���W�B�<mk�H�K�fs1��]%�=c�6a.�P���������p*��_�!��n�j��A�oS�	���a47+yH����N���w)�m�Fh��f�Π��.t��i���9�0"�'�C-6���$���,��0�0�m�0e��}_��t�^�+����\�?�%v�<^t��˷_�j��8AdG�n���mL�[�$UKY�LV����PN���{�f= '#^�wgoٰ�@W.
d�H����i?f����|����x���|�I)�e�Hˁ�M\��#E[!��cU5j2�y*���|�^���4��?��I�!!ح��q�Fb5u����cA;�Z>���unx��Ii-6��#����[��z{F�Z���̅��W-Y���تiP�����B ȵ'�P@�M��~�An���$c�U ˸ٝea��0�r�� �t��:�n �����Q���U�)��%vrk�͐���/�XT1�>h��p���b��k�^�w(�$�'�Y���i6�jvM}����Qs��so��&{�7li���n�R�
�(��٘D�b���K�|z&�@�\7�j�g�dv�����:���骼�Y���R~�ڃ`u~���C���A���$$��|0l.�#$���l�O�>|;�,���|��<NQ�����LBP8���K��* o�*�%�g�,J�V�b�1[�o�_�T^�:�<�W̬�8�I��mb��u)#���&��!q$�>�Ͳ)m�}��e,Lmܐ���YU`���6��$��'��f�X0�e��k���e�6f���P�M�E�eX�sǙ�P��8M�)d7إ�ͱHa ��������a6~���ܢɇ�c����!a7�E��p�ՖΚ�dZUˊ���o�B:����?��酋��j�"��<�_�С�]F���~��$�ӗK�x3��˜j<�?���Cv˿�WQ���e��)6u�̄=i��/�Y�&&h|M6��G�<o�&���g�Q<�+Yi/2Zo`	��D��I��'H��+y+&�
�Ġ~!���^vF�Yh�,����[<����d�$'I�]�A�&*�F��ZX/���`�<�o��	�(V����CmI!��T���f?��D#�c^B�)&��B[^a��?�K^� ]�������T�scm`f����ۜ.a������Af� r<?nN�E�o��3ĉ<�[�֥`�<�_cB����c�!W][���*)=���CeK��ֵp��h�#�?�}��\�ߍ�x�l/��;��g5��O?�Y�gz��\���eX$���6`ao��~7w.L6-V�z��|�L��3�?A\v����؃X-�4�������Blc��RK
��.m���Ep�p���"��$q5�"�0�fN�CET�F�敹���QJxR�r��2�����Ëg�������ӽ�Q�J�kK�Z�(`a5]�3"Zg�����9�0wa,��)pj>���1z��pm���Ҳ����L��M�O`�{���w� T� h��U���_���cdd˟|�"%��KK�`�I�q��P�������LO�w�zՌ�\�B��FΟ�(�~K+tB����}��]+6}�:�6>�\!^��M��b��s�'�q�pO/)�����Q1��ED_��Y"0�iIQTOZ�Վ׉Jh9Sq_�7�nq����[B�<��8�۹��ѽТ�,�@��s�n������o3q���-��O$Y��,v#����t>�YȚ��� l��� ����W,
\��p��O�A	�]ᡑ�G����E)	��:���=�N���ӳ��)6��NGd+�����Yz�ܨ`]���d~E�Q��o蟄������#�X]����EiŌ�(�QE�g�?G��w�����P{����۟�y�f��n��ȓ��-�:u��,$�����)7������S��D�/V���	A]/����Bi���˅�d?�<�k�d*O*�F�~�<7�����
�t������6
����}�\�#��b�_����,S�L]{֎E�oz(*�2Q�]}� �nx��}lƉl�����E�'6�vӯ��SG����M���٢M�����y�ߴ A��r�yg'������\�t���k����˺�dF7'kJ��F\<�s�Sے�5�"n���g�z]
��I���HG7V����6Ȁ�\&�?u�m�"xNn�&l��~�x6,��yuÔK�6T�d����Ŭ����{�Q��*�eN�Dv.��㖌p������ȉ��m،����w��sLq���:S��nO=1?�җ
���`��=�dh��a�NT�R$���!�ėq�=���l�~(u�L�w���=�4Y�X_���f��L,�����&r1ۋ�aά�����@L��ߌ��Eھ�Jkө�ڲ�I ��.	#�8�l�/�L�V	0��v�v�1��M��~5\�"U�/�F�����>���J�UɲZ��{�P,�1ԉb��> ��/ e��9��n��:�U%=����9��Wm
����ң�8;N����4g��O�-���tv����+��|j=�߆: ��gTއ��p\�{�R�,r����̖��iۜ��䷊jm����q�e�q�ΰ0�4�1(���kr��L]�m�er���A��_<���ː����Q���@(D]>��3kQ����l%��v�7��c�GWm�f�s��8����q���?�=�5"�=EP14�q�3��8*���`ds�U����S���6i��5:����˄ ��4M����1ĆNJ^N��*�Q�sg�q*�y�,����ԍ�WԀ��8�B&�D$S'z=�'+�@b�.:$�$�0���3���G�:ک(1񑸕k�!�^�ņtnxnз��@�T���9���A�JbϏKC�C�܊�>v���aN�'m�ю�^M�ug�P�p����!Y) S��t�B\��!=�~�LJE�d���c+r�%��s�G�؂1�8�G$�(2z���!jƶ$�'0FRh�}m>���v%L�������� �k�O)�A+��Iِ�.Uo���a����dQ�薬��ң�BI�`�������[l��M�y~a�t%��m�U{쉺��<e�	�l�����LfIf������3�WZ��y�X0HR�eJC�3������n�ʐ��-���E��8|)��'�:�L���ˊ����«��!cZ������(��?ɘ�7Hp�h��Ә�=<}�oG7=|��K���J�	I��D���c}�����)-����ǡv�(B�^�#�R��"忎�c�Z.t�����V����0SۜK0�d�v�2�l���9��-�ؼ�"�ɤ�[�sZe��:�P�>�P�ʤ�Y!��]d	�f��f����ū@���˜7�f�a�]�Zo ���E�(<�U���Vz4�:��a���L����5D4�R�V��,B
$��^�l�|�zZ�m�����Y���zO�`�&�>?(C�2O��`�_�s���r�.�J�zΒ�͘s�!��t����1�9���2�E��Ҭ���]��T���gU>���wo�-2:���-C��d�Z4��#+��$����!�B!�,�R��},rL+�uO٨Q��ҽ|d|�/<H�芀�L�e�B�ɧu�B���L�qw�Wc[�D����5DC+u<�M�)1���b1:��w�c���`���/bi9�Aa���Y������x�z���<�v/�Ё^���ѿhzdV��f��h��B e!;{�d��}=�[񤭝���'#�{��uI(y�(�}/������F�C��Y����S��1��o�G��Q����c+��D�sB��鏡����<(.���}�~ �NN��a�դ�������Eg,Q�^��	ѩ�f8�~?�G&,��mS�]{�g%�0�)q�������L-|��@����,jy�5�@���T`�ߺ듙��؟���.i(�̵�'a�����s\˜��h�/��s�z�j��E�/_Hꈹ.WZDQ4�v�Rq��b�=/��ʁH�21�Y��ȗ0S�hu��H����n����i%mU��eu��}���3�y���'��
���� Wg�ҭ���W�>r}F�\&�P@>�N���0B��� ����h��.���b�rw8��	
ZS.�o�������S�r��z���p��&�t��q�|X�i-ٕ�d�*�������E~-��뉼�.lNe �2m�"��8Y�i����6�Yi�m,K�h̒���2C�@cM3��.ڷ{،�b�[�n��軡����R�w�Dy�9�}7��9h�Gv�M�f�!y.p�LN�/�_})]�
m��j�����r~R1KzC��A}Hp���B�Dd~-� )���o���u4����%�w��7T1�WG�ؽ%D���<��m��`��i�mT=�����jx���Q�<a9���#�&Ɍ|��8na<�3w�!��-�@�O�O�#���Б7�<=�%��GG<��O����,�ɵN,r�&[f��Y�OD�t�,׻'^���������O��BD���5��}����h���5���@�����z:���G���Y=�.Y�_� ���L0z}���LS&�ꫠ��j�n0�����\lR����~$�/�R��1��������?��m���+�R��l�c��g��偗8���c���S��A �dCw@�cFd�z��!��9W�K���0����RK4"[�\��`��AY�Q���|�*���Zo.���3�����d�ZY��nj1m�1�ćyv�����3-�2<�3����pĢO��u?2Թ�sջ�zC�(��$�Qz���%;ѧ:��:US4���3���/����9Z�'�	���_�,l�w��A����
`Dh���:��9��D$��s�9dw��_t}��m��e�sKt�N&l�B��k����o�D!�"�>��}_�;6�1x�B V����@�m�9%��ʫ��	xƋIZ(�i?I�}/�(W����u����J�����z�[.�s7�7g�����'�4��t@)y3(Y6˶cS��b����Q���� J��5�����]�Jfj�3z5����$�l�r(<�׎r�<�
����C9Ȳ��hF�wW��{�6�6%���q(%�,�t$��9_��)b�p�,�r/�̳�.<�T`�o�Q�H��;E?��
��w�R�Xʷ���PAnnQ�>��{��6�z�쑅�ˈI�ݷ�/���P[!q4�^�/,Ȼ�H���w�W��U�^o5�t-���cl���F���ǐ�WN�,!��,���;�.������b~�K��eV���Sǋ���e�!����5QI �qn�c]G_��cd��Ǣ���%�ݳ�+���5�N�bS9n�vTE.��:��w��kl?����yK��q`�6���E=4+&"���*Y}Ҿ^e��7 �tX�Cx����,�e�p.���q��d�7�(S���ͭӬ��S�Zj���o���|F�a{���Rv���S��ٞ��:5�Yd�����~?숴��Ae<e-���&=�x�=|O�0��G�A�+���73̟~�
�s�:S�D~o��1H��G�7��F��L������M��6a�θ���ew?<�ҩ�>��HA��Q�M�%�i�P�#Vn�z����:0Be�MOو��ggꅏc�����G�:PLA�6k���2̖$�\ͦ���0@U�G�˅��u���b�n��1��-V���_ŽA��#Ü������sh�)�p�g�3�7��Kݚe �x��2P�u�͖d�E����aO�X�mGB1�Zz�MlJ$��
?�\F�B�S�҉��
S��~�nu�MS��~`���7JI��,�fO�����
�c����-pD����T��܂{�j4�7��S�A���S�&�T��*%���\ޔ�[����tau�bzJ�D{�*'�w�gȒa���¬�5m���AA�*3��m>O*��-7�m��������'�y���.-p�g!Kh�J��l^�?nJ�$Xb)�r�R��}���7���R�hO�*�#�&������t.� f�t���.7��	G�g�{Y[�^��
�L1�[�R�]�r᫑�Y�Ye���ÇތN�c�ҺxU�N������*���;K�}�O?M�#�c������.)�a��Y�g�e�
a��4�O���n���H>�Gv6vy龰�e�\|�겕��?��u��5;Bق����i�UaWv
�,�w.~�W�D���`��t'r{��N��}ķr�}Ĥ�|�&>,����r��&%�85ϪO�I�loc�#;��=7��s\�C�x�/��r����_]'��R�'��}��=1����9ѝby���޾�x�]�?�8���<�}��Շ�m[�̿���U>�����*0M��y>^����(�Sn��B�|9E�F6��oK_��xtJz�k���8�&>����Zy�
q�r�*X��.&���{��~�,���Hd'\�گY��A&�nC �(iFU�8�*ƌ�ˁ���.ᭂ�*����lo�̊YNs�z����m��r�B�5!DӅ!�\����Z'�ml��i8���x��,�����{�����B���H���m���6�ƴ�8y|)�Mq��i,���j*iP��҉���]�<m{dL�r�(�;���A��E���1>��Ġ��K��$O�ؕB}��1(���2����ݯ|�u���v�P��.w�W���{4 ,ZByYL'�)��Ԫ4w��{��)Z���*��m!����W����
xWz1�7��|30�e�y�1�3:�Z�"�R��j*ź���^�U�u5P�Ԙ�tE۽�:���ղe>[=KR9��r�T��S�N<KC�m\C���]~�d�B�JG���g	�����e~��k���bAZ�Ŝ?f�Z�YN.y�8����:Ϟ�0:��|���vE�>��I:�$V���ԥy��!����1_��ЧQ�"K�Ԡ3qM�۞�*��m῟���_��䥉�2r��SJ�������mp���b��ؓjI{$r���g�⥡y�t�z��)v��ۼգ�i7��ۢN�����ry�;pgM(�c�]�X�lF2���=��,�D�`��6rd���n@B@t�æߨi)\_Ԏ\���E��*��σ�ҶA��ߚi���G��go��\;N	�u���K��s��x���x �p�/[U�~>����Fh-�c�.��Bg�\��*0�������6������R	��\���Pm�^��xO��y��P��-H��+�1��8fӰ���$V[&��m��q�iq�(�ڌ�0

�GV9~��_9,;#��jٍ�w݀�������u��V�sk�Lr7]F�V5nT��:��
FW������v�5<��0nTz�H��X�&��U7g�Ĺ�O:���n�QY�dJ�DB~�4U���3����e����������2���D�r��J!�5>�8�����Cs�w�ڽK�Գ{���+/���Q�� ��LFx�e\��{~E2����t���-�@��P�>/(�Q^��)ڍ�xm�VRe� ��@���*�d���7_	?��irpZ�p"�*�}��ve���ž�Ǫ�4&N��8<�w�M/�ꤿ ~�,�i����|�`.5̙x
��YI���/_'��Fv������$L��ә?��4�r�Y�yz��[����`l�G��m�/�1����'�Ӏ����1��,ϔg	��wت�GD�T�t��ixF��$i�o2P��R��bg y��C�n�2l�j���� \JTᗇ��}(��|SM_D���g1��cF뭲�o����n�o@[�_)��]>w�нqN�j���L�ЫSS6�U^L통L�s�>>Aw 2��mA9X�[Y���/�A�E�f�8HC�i�&kW���&i��<w�0���y,ax'*�ge��[X�b��;��LD�v��l����Nn�[��N+�k*#/�~�|�U�A�����t�3��\��hKe�#>w?�3��< \��i2�8�&�r6�ghθ�U�a���KgzT�McGBl@���Df9��-�׬v�Z���e�H$��hP&��+}�&Z-4����m�0��3Fc{i�}�v6�V{�b���X�Ӗ���6Ӂ=�o��f�6^}���h)���%#�<��xǾ��9������U�#"��.����5�9j�0y4��t��M��Ke��m����V���a\�@�㊨Ӄ�V40BT��T�m:�ۇ�MFE�D� gq�>��5nn��WBͼ0CO.�c��}b��Т:V�Z�N]ܭ�c���_���*���߽��|J�R�%l�9�q�
�4��n:�V�������S�ll�׍��ag���f�a�^4v���/u�;�B�̓2�S#B$���*+2�w<�6���Q�^�V�n����5}lJ%�_����ױV��L�sz�$�M>�|�?��o���n\��O�3�W2=ԙ�K8c;�M�������7aQ$5�����kt�O#���v5<��F�m��ט��8v~�r9nE_�0�-����؂e:o�sF�o��'��	��AI�6�e�$�u��n%Ѻ�k-�dOQ�>�.}/U��*YmOD�!6���P����JH� �Ǵ�H��3^(��X"�pF:���-�H�#�VE5>:י�q:����0��d�'�����go~�}6��Px��0<~sQި��c�m�����Q9@�z�7ۦ��̎��-��oqo��}� _��s�ݘV�ɢz���s�����DU����(�^Ո�ꏓ�����(\o�t@q��Ñ����7���xH
��}�FKXG��^DGFk����f��)QP����$උ߼����͕nuw
9��Pv�	u�R(��l���Us!M �b8����x$V�(N�;�nӹ�ݨ�a[nG�.K�����>jy�X�"���\^umA\��)%�,�ۛG0a�L�I�Пxb/��F]�]���)�"��1�CM�^�Z���3lyC䷳|��P��̞W�ܵ�;[�Y�p���^�^',����R���۬���J\��E�x�t�`Ժ-�5$P{D=�w��
�ۡ�y=S�����K`��XU�	�@���h�XT��(�h��#��ږ(GR�x8ʟS�������KX��|�tH�3�-cd� -Ӽ�qd�1���L�~Q掿�ٶ�]X�#����Կ�V�9���`]�C��Ю��u�Ч��o��C� �R�Қ��?�I��_�l��
��9�~\��2��Oy|�c`=.�t��2���ӿ�iFJ
�_��4�;=��ωp�_������BI7r���S�o�$|l�4�����l����H��{��7kqsZkF�bK�+~r�l;Bo$��C�K	��9K����*�|�}>�>TbD�)�*�R�d�4��ٖ:8/I��.����m�����f�B�TDg]�p��]p
0�%�ݞ�(XQ�3���w�S�m�� s%��ѕnCp�Q�k������Vڛ�X�_E�#O\���:�d�9�U�4�5AIz_uC���4v�7(OpR��۬�����@?d$i�I?��AX�m� �wE[��f�-)�9��?�ʌ���>կ���B��j`F��r�O��N�u�-h��;z�e�}�BLU]��[b������������1H2K��E�ܫͳ��
�/�����K��șg(��H�C�JLQЊ9��8���.�_+���lvђ�X��mY�Bz��$�(��Kyl�o歩0C��V�޹z�N��f#���C�`��Z�'�`��[�z2�J㐺NL�����=�7�M�􆘒��1^d���HK^�e�,=!��l_G&�|�����Vu�Z�P �����@�����s+.5�A:xl �<����{Z�~n��	��1M��?�ɩ��ӛf�������nI�*�`˗�ƻ9��O�����&�P����
�؉��0Nn����	{H�/���Ϝ���CI�tDoz��aI���+�Q�i��m�m���n���H���Te�MP=NtѤ�x����vU�O!�D݌3$s���))��	 *;��� '������w
On����\�-�V1��]/�w�O�A:rb÷p��"�!ВY>@En&/�:�8���[�i5�,?O�h����K'�N��7���s �{��m��uc�3���2��9��/4��e�N��6���S �ET�/�N9l�*���mY$}Xo�����Q���/u��9q&S�%��"�� mC�!�{��%�YF����<W�ہ�͑3]���Q������ŉ������uΤ?w�y@�|�;?�c����u�h�i�U�%\q�>���Y!gA����!�͏���n ����*mfu눖����m�3�p��4z�JDg��$�F!@��c�>�٣�P�����A1�D�>��>��t,US��!�[h7E�VZ>� 0U�ՓE'���{�x����������c�#s�E��:'(�+1r6����;����ɀgQ)D-���9`*���M�kð>��Џ��0�]'g�#�a���MnN��S?���,�B!��s�s��R�^=\�W/��� 4/���a���MY�̐���񠟧N�}��N4O���XQP��t�w@�{�@�g��X�����Q�gTiAU���� ¼(��K ��z��@mq�T��s��%�UZ�1�����B�a�@�6�GJIn�>�eZ�V�{���L\|�U� ���#S4���L�z���p}(��2�:�\	��ٍ��H�5bI?������|��5{���^�pT��m%�1_fŞP֜�k�6��r���5)oLf*�IZnE�H
�]^wnm=�T�J���S��`����M��͔Cs���l0��g���>+��؃���}���]n�X����<�.&�����*�(Z��5ʕo��p�
����v�-��W�dK@�7��2�����f���������<��d%���J�_��蹾���ҍƟ��U������h������K��Z����}��3�oضVB��ŗ|[i��?�.���/��c�ŋ����NY��Ɛ�	�^O6v��ҋN�o����W���	~[!������_bs�J��پص;$RbZ�y���eG��U�{���{�6�j�H��+`B��m��4r:���Q�)�9���0��>��WɆԣfP�~|#q3��쮗���3�I����'��bu���b��G��L��6�,�Vx����v��67ZL|�Wwr�
�o�+V%465^�_����y�U�s�k�'�F�����Ő�U���b+���|�o���>�����1�G��l��c�~!P�
.��ަ]����>=|Z���}�8��Ix��@j_{���#)]v63��|�[X���Y�e��>گ& N�0̾x7#�����(�w��fy��[ؖ�+�s~&y��<�{#ۜτ�+�e�aG6%\BK�C�J�ᦤ��'5"=7i*}�h��'ǀ�A���og�ږ�w�c{tI���<�hl܌��M<�o�������KoX�n�����P��%��N�pjA����ֿOZ��8�1g�C�;$�vK8Ka<m5����#���:$"'3b��)s��l��s�$���]�Z����|a|�C��ԌW;R�z��y�����{��
`P���hRVys�q�驞�Ѻ%x����4������l�"���X���cz��[�,ޞ�j&�}oZ���^P�zڥ�D��#:^�2���[�c����2}Z>+�C��p��]˄�
���/�F��5�f�g�pWtᗇ5!�5���%i/�f��4�G��d�(S�����¾,�*��@F�~J(b�O���r�*� ����a'�J�����a��u�K�A�{)���X���m�V�i�K�j��aX�w�h�H�J�֖/�uuΧ��n��0
��bFEZ�e�t�I1�W�u���3D�����f����"�FD��c
$�����D��C��zeEz�#͉y���,�3ח�ܼ.`/��Q4&]���ܒ���V��~�C,�Y!J�W�m>�\�c'I:H�^�E��ʙ������8�?�*������v��];�N�5<bI���Z�ĉ�Џ5ʁd��u�4y~�5���ef�������pt�n����ܭr٨`a�1���}��B��b�ڞ(�Z�{�[��|�7�֭wT�U�_�"������p��l	������}-Nɉ�����MK>��'V�|��I����24�7V�d*�� ��ŤO�`�d��k���1	���	4�C�E	�>� Ⰲ�y���D�L�D䰘�(_�_��ZñU���}��̈in?Vt��ڎ�BfU��U�H`jԺk�1T R�>iD��@@�ϰ�|'lf�E��u﯋P����rz��f��S��ѥ|���!���OϠ�{��c�T����i�R����$@y��2G�0�	���rB�>a�+cF®gAn��'�M*�^��Sݻ����G{Q�yL����Z&��hD�so���p�����t�$:�	���:Q�2�N,F�׻�����g��A�3U�3��iz�ge/O~����-��-	d�Y����P˾dG��f�"�ֳ�a/�7
�{=j�\���v�1���^Y��r���ˎR�@|u0OzQζ��!��16A����U��6�N��0��}�!kX������Dh[~)J":zU(z ��թ$i���������Ӻ���^��4v���i�j��'���@����b�����س���8�y�q���<���'L��9\�\���<px�%�(0��#{��z�֘�o6♤���̑H0�w�>b�T�r/ukְ�B@��h�U7��XC��e�W��� �+�Ei��9v�zZ�C��o=����Dqp~<�W����4,��4��z<��W���B*���\4�V�4S����?[ϴ�A�����v����[#5���HzР�{��?�YW�@�*B�m6���QG���=Ƥ�����*�m�@B�|���wx�\Cgk}A����_��=�y�$�-�YT���%��$Yj�%F�+�{��][j��W~i�G�cQ>�,I����v�wݕ{�rfz����_�ǡ��J�7��Я��gnM�W�_#J	ǳ��މ�aA�y˱o�9�jfN)~��'?9��-T�4aY
jꥨA\O�=�$�:�j�H�TA�89W4�t�tu�d�lP�{̢����|�7�Zzy^�9Ϸ��߭P.k17��T��P|N�l6�ގ�|7�=���|1�G�rX�!����b��%�%�c�S�^\��=ub�ѐ74�����}|FfGy]�U�� �w�!�_���>��0/䱪G� g��R�_����O�D�0��ߘ��S^�O�شVL�ңh�k�˨ާtt���j�Ɏ�� �{�d��f=�,�t�����fd�;{�M�|ǣs�����E�G��� ��r7&0���r'�Ѭ3�,��w𣖯�t]�����W%2p���70YDv��U3hYp8	!�4�jP���b�[���ω�NÊ6��2!���"&8wy�S2��QB0^��lp����_|�x���WR�m/ʷ򞍢Pg�<J[z���D�_ �q�%�;z����N>�Q���ν=cQk�Y�K����Ƃ�q�=�ꪭ��v�qq~}}}�X8������?���J�qu��2��U���䢥ԩJ�'��I7#�ۏe�<q�ʁk�;eׁ���Z�Nܸ�<���}�p��{4�;z�gT}n�!Ѯ�W�dY'�A_�[梼�[��]��k����G�\BR�Nv�
]b�c�sG�����f�IѲ=���N�����٩���ۊfY�T1e��C���A���w'�7�����*˔!s/x炳�����0�ח�o��Ũ��R*d�?u����):�����v�'��p��������E�=!�'��R�Ml���h�����������~�73
e��faa���~0|N[|�M�@B,���д)�FF�������K~>��_���ݤ�K�i�3��R��!rA��=�&Z�	t�U�Ċ�U�]��bM9�T��Ql=dw��fݢ�c����A���0�km���W��
)��}
^�tQ	D��;793�H����%-��H)��e��F苋#Tqٺ����&�w���w��{�O�Dx}b"/�����@8���Ǩ�ʵ����Ƴ��=@}��)��̊��}�5�Ϫ�i�5E(��V:N~�5\͟El2��i�׸��Ls%�[���GQ}bB����<}$O�Rן�\�3	��
cSy������U��n�=A^�Jg!e[�C,-i�E�b'�o���e���O=���י�9{��9�{����m�YI�哾��@b��pn��&��B
[$�f<��O*c$�/�ɍ\*��1�� �ׁ�6��=Nt�(O��qrt�#���<���X����������&ߌ�ʼ�I�oy��Ϝ��x��~�[�A��- ʇh�̸���]��^�8�+@�ߥ���^%��*�]~�{��L�vݨd<���ZMĔ�.�lU����$����TG��&c/��/�,{�ݮ�����XA���|Gh���DF]Q�SI����Mf�e��J�j�R>y2�D����!Kz[���61r��V��k��ĝtg�\w1��۟�})�U���պw%h�?G���J������͏m��'���?�ug%������d�1���f�Ӧ�����
8m�J<��7[3Eb<S~Q��X��<���jz�n��2��rƵ����ư$݂��+Fу����3ʤ� ��1�Q㦳>��+���/T�,��t�grf]���m+��ͷ� r��gX�_��Y0t/G�s�k���}ݺ�����o�����U���&7()��2_�8��!�Q@��EogL:��n��?
�9�a�a��1]���!��<��ޔ�v!����!�6��L�l��Lۄ��׭�;�L�?T^]�9\sI���|�������e�l���AM�ɛȋ�W%���B$��i������8.:�3�s*�r��o�KaS��s?��2͈��etȝDRn��،��nnm1�n46l�ݗ�7|?�}~y}^����z=>0��ݐ$~�p���[��
�0ľƓ*/#.��H�f���K��\�����0��s��Sijh���, p�C�(��4b���tbh��e�(�)N���h0!`ꯉ���@�#�-�dB�k�>��MY��TY>��3b�^���P�hw��h�&n1�k���a7h��u�����z��,�:g��>	{��-r�E�?9Bu�h�(}I<��D��r�Wʪk�7�?���ʈ�6"�s��vӪ�8��[���,�"���7�)Q����u�^� �Lc�ז�9���z5�An�%)xcf�z����c��*��� ��x�`?{��?$��F����Hht½��Bԓ=�%G �ݘ������e�C��S�	L-�p���(�ut�89����Ɨ0��U�� Wl��|��l�DG	R5��>b�D*�S��}Oଇ_�zj����K��9�:?�d�D��<��{��ڼ��"em�I*i�+Pź叄s�]���*4
��^F3dʆA%���;��K篜>LkHJ�Pw�Z�f�u����7�-���
fQ�>:J��D�|�u\h�dН� �ގ56/�h��g�<o�$�����+��A	��J��L�*�+*��"��44���I�v��;:�u������(X���1}.[g��X�HR���a��R����ug��7>����?���)8Ef�����ҞbH�d޳Ǌiҡ5��!��}�[*�7��]Yn�dx~e1R�O�GƲ=/��\M�9U�5���F}��݁��D<mWz椷�J����\���iA�������k���uQU�azǲ�t]�~��s�S`��ځ���U�z�_��U�I�,������ьyG�'�0n>O��Y�!g�;�GڥCjnX]�Ira�zh�� b�����]��wð)<�8�v(��o�C0��9��߫����*����tXk.&�W9��ѹ�7������u�R�N����f~8�E��?P槳���5����oٰ�\&'�K��m����+O���8��[��aG̫f5����߷g~���ҹ.K��������A�y�y���+���8�N[x}����q��û�N�+����YJZ�;��=Jް(�E�LXpߝ�W�%�������\L\F�UM���#S8�A����zf�\E�E^/��v�l��>t�~��k�D
qL���s`$��=6��p�*}<D�����9���qͫP�M�u���M����	}<[�ᵠ$�Մ�%t���[$'K��}�`TA}	M�P�3v��5R���f>V��(>��'��R[[Y�<q9�����[|��1��`���/�|<�uCw)͛:����(%�ػ
�=B#�O_^�܁@>�>���9���SR�B���<[8�z�MQ��)�K���nD(lJaH�u��q�Ҭ�K[��[�k�7������2�m5�{lm;��-�vȖ!4�yPs�Kl�ܱm�)�cDs)}@���U��Ѧ�����0�i˗�9La9����/�����m����`����7����7����3C�@6R�HR��Tp�F~Vi�_��i��,_�PB�p�'�)����.�#5��m��vv<�Jw��.#Y�4V�_鐒���r�k���j�X���(��Di~�@a7!A	��?��kS����T�Za�Y��G�i�S����#|D���Aﲳ���,<)m�V�m�b�q�BfI���'^,�*� ����O�"�zbW��0�&T��vQD����֔�K�d"�֒�{�R'������v_�H��>�}+�Hù�Ė$�#"�'����<Zw2��q�����,b���.3�k��\VW��-�q�|�ɯ��]���\��5�j�j���,z
��$��8^��m�ߜ>�酳Eu�&��7H�e���ډ�QO���|�:�f޴*6���վ�8x2�+�%�0�ˌ8�ˆҒ��j�u���_��,>J��t��S�Y%���E|�C�Я����� 2aoj�ꫝ���?>9�.�:l��-�f��9
��v2��<}��[�b��@��A�x��T����������-^����	�!����iy�p��rU����5Q_}ĩq4@��ܥ�2��i_S�ƽM�7\=ń��=�+��:{��5^|�C�`�5�l���@�ye���{�D�@U�)<wYJ�����1rh��f`�6�B�oX��6ǹq��y��6M�Y��&�cSl+{��pF��՟Z.�V8$�U�xn;�ǻYʷe}
�Q���ܱ�.�秙���3s��S�%m��Xm�vĐ�������9ݏ��f�rlE�+/�\��*@]�<B�Q���e���H���m�2��M��1�\ۮx�sXtܩ"v���Y,!���Ok�r{]9�������:�3��a�[vyau����٫���y39�{�ώ$��|"y��l0SFH��]���O_S%;A>��"w�#�z���K��l��[ZaT�zOC�؜�a��T
�z�m<�˔gT�� }�ty��T#A�q #�V:�w�0)�b��˗i*t<{*����1	�<�;��m �>K�:���!�¼����T���V�U�U�p�j:��Z,���B�%�<@]~��M*%�3s�X�{��;~O̬d���|����0n���XA���O���
���^W����k����X��O#6Aow^�4U ��~���P����T6���������;�g�W�(��h�=3�#>��#�nҨFO�T��8����qT��7PK����.��2���\��`�ݢ�]s�!�j���߃�5�S�>��Z���?JܔAIB�%���&��!�(��j�Z�wCnT(U�2J��t��+���>�h�+{��y��_�X
ɺݿ���XS�Qc�0,w�cN@􁩭�'�g��3B����+W����,�S�n|l�^��(�}��kA^ʊؤ�Ԟ�!	2�o��f��擷p����
WxO��c"��@��<�h�,�(98P;K�������at�;�ޔ��p�S���âm�/�#k��ѠYh=�e+<h+W^y<�/����V`x9Ę�s�M:֕u��h�	/m���'��s�,OO�"߱���$g)=U��)-ieK_w�T!�d��pO��\ɻ��g�5� Ht򚶵�E�#U���9����]�G]��|7�^bZ[���'�v:lJ3���e@{�	T ���Ȉ����,��m�[�m��*M0ԨM�W�(i�
��\��J��SF��}��.ڄAu�+��l!�#`���
�.`G��+�].R{`v�m~�S��|����숽 �;�\��.F6�T�Q�1{�^��&&Y�WG��9�AT'_�HA��B[NX2��Gޅc[j�U?��W8��F�{Ŝ������L4��?����o#Rh?���)�Lݪ�3�9"�mR\�6��A�:ė��Q.����Cw��⢸ƕ7�صzʋɄ�\>��j���>�@J\�6�t�n�Z��K>y���g��~1-�w�빼Gv&��7�<�o�/
��ছ E+�eO6Ug�b�o�T��T�A���c�?��Y���;��U�J���v�b��p��6��������3،��-8���Z�b�d��@��?��S�#A/���H�EE��Y����5�B�7B�x��w� �(��q�PK   L��T���"d. -y /   images/4b94d0a1-8bca-4ba2-81d1-ddf4f146611c.jpg�}	<�]��=$%�J厐��l�X�g/KLd�+����d��!
�DT�T��"*BF�5$�����<���������{��O���9�:׹�u��|Ϲg�=�f�®����`0d7\��G_UO{;��B���"�1��!��`#����\��0�{>~x˼�8�]
�-`	�������7;��f�*�́s�DoI�ACW
��K�o��:���k����K�%$	1	1Y1IY1)^����e%Đ���s^��J�||+��j�F�E�IH�3��y�t��wCsqNC�:�e��]g>nq��9��^����d>��>����3#_<��a�3ȭ���� >w�8�<笠�&���cH��1%��87�8�|�8�Ť���OqƟ�R�|���?ɗ���V����R�S�Om����K������S��V��;�E?jCy�k���f^�l�纀��R�1�̳]��E�8��5,�?C~��+°<�C6���� v"�z�NLO��,><�����֎�K��Z��ٖ�L�f��o	������54�#Ǿ�������?���
Q0)���6��C����|x�oU��g~Nj���Nkb`Pa� �3<���Q~qmXS$�Aꀋ ���2��a`�bipS��8x� %�� ��.({�9k������A" �#���pGC^<�C=���� ���'����Ѐ����@�J��:'/"H����������,q�]���r�`�.�K"�C�ȓV��A��W=UUU���T9�#�9U�V�[��V<�% �)"�u���ΏRn�l���{��|w�̃x�e�D������z�Ho�?| � �N�Ύ�y2}��Ős���k��B�
!�!��lJ^K&�$��]�dr;ٞ��)�������l�)���L����!�%KA�������F>F.';�c��dOr���'������cd2�(9��䛠�\K~XQM>L~A&�mɑ����q�Vr���L~r�jȋiY4]�FH��\q�}4àdY����o8{i���c1Z���ˌ���Vz�ќF�q7៺i��tj��~�5^�7'{=^2A�qm�������������?��'��G�R�v0!o���f���7��	z����y��4�x�iA� ��F�ͻs��]������1���~�/���ܱz������Z��׬��fO��A����=�~W�������4����ZX��b9�O2��v%V�V^�L��UYR��P��Xg����?���t%V�}t�>]�?�t��TCL`��k�8���ìcC�g�t�\�{��zH+0�l��n���0/��Vt.��	g��)��IgsTU�4��8� ����v�Wo��7h��3�?�-T��_��o��۬��a�W����6���М:�T���MYh;�k?} `#ρ0�X�=A��sO�f����p�~�_"{����DZ�����.{H%�;W� �|����)�"��@x���hnG�ѿ���.�Co�Clls+%4����Ր��jE͡S���T*5�z�jN=I�C�I� ��sNQM�TG�D�J-�
R�S�B�e*;��Rc�;���k����:�#X��
Qc�7�Y��>�5�:D�:}�j��ğ��z��@���P�Q�S۠�Z����L}��|�8��$Q�f/9�\�j����n5f�]�����a�W� \��\ 4�cY?l�`_��Al=�d$	y,� |O`~ >�� �q.�=(�����j�6U@���@O� \�A�mA���(sYu���x!�X'�<x� WN"��bɃPJA(�$�A�a�i��@&zK� ώ g��o��� js>����8Z6#�/����6��nx6���KЯ?� �Y�C� Mɀ��_� G@Wt������������'��o zBf����t��2A����x	��P���L�'�L�0���"��45�)Y�p>���Π�b��*���**Y��=@_H��$
�}Љ������덦���h�=��E��׍�D�)�--�&\���"���9�a��NÍ��~�S��a��E��1� M�ЊH��D!��>�r,�/~�kfF����;}a����9`%�O4�������N����U��� �i�Ї����r���y�LA�6�E�5P2�UYP�p�?Q���x������՘�i	Ӵ��t��4�����šj����ܥ����BXA{`�A[Nd@���|�ZM�F��a��tQ%}������8�%��h�R�iZ&��������x���h��#.Eˡ<!
��/����V� V@�&P-	�K�ы�&�=6k�>��ɛ�A��P�r��&���Hp�,Pe�Ǡ����4��"��6�Ȅ
������ �_�6��D"��0��ɥ���W{���@+!vCY_���i�!�=1&FA|�.|�=$$��[i�<���a�6�k$���z�EЇ��EX~���s�!��#~�I����w�� ���Km�-��X�۩��Tw@��k�#X��cvQ� �R�?R���#���g�F�i���9]�K Ӂu�����Ϩ���Klf���E�,cL�4;�!��1�H��2���zV��I��3��;@IY�E��J}Vn���Գ&�&/L>�?����%P_"�R4,\o g��v��u�e��[���� ���ͥ����u���~���s�����/��Mп�Oʰ�� �@��N�
�0�u�����L)��]�[z#�g�up���z� c�:,A�� �7|?�էc"��. �{w���P�zW�-D(�6ؠ�J�S�{�y��zgu�~��-� ��n(p+`i	�C2 _��*�t�}��&���l��|Х@��6��kg �x�#��٩� ���$��B�5�}����������%����.u?�K\�.!�K��t�����}�<8���sl>p�!�y<�K��Kf�m�����n,�/~�kfF�����n���a�_�����Os���E���?Ǣc.��/ �JQD����Ve�т Zk ��qg�g10τ�`K��v�O����?����h�U���2bi�_����/ХWQ�\�^A��b�mS3�#ڧ�-��Z�,�@ujS��	.F/(��K){kjP}��9�9m��警M:ь\mʍ�m���@5?LQ2��TE|F7�z�L#�#���P)	E�z�	J|�ʶ�%����*q�΍��e�Fv6���g�7��)'q픰�8ؕ���vCx�F3�B���H�Bɀkr]�#�@"��q�bZÏ�JĠ�$��\2�h� �*��ܯ�\v4�J�@-%|�R	,�m�$Z_�F0��5E�p�%�t�s=P�\Y��D�+��*�\�K(.��X�3�s�F(m.�S��\�>�D�rQDb)%�f��=����>��"�+k�P���.m)�`���� .9Sը����
�O�A�� D-���R���=`�#`�`��AV�Ӏ5}pr��8����!�)cT�G��Rw�+NB�p�!"��ۀK+��*@�kp
�ƃ�]ԯԽp^��y������jk��D�(����<Y��!���>��5��+�,BBa=���=�B8OA��Q�A[���u�KX�Su ;7�C�w�L��=�A����P�Ɇ�a�%� #�b���('�&
:!Ā�%�?�����nON��
�
���؛��7Ƴ	�vv�A�c)����pO� ����Ґ~XE�*`2���P ����A���·����� z����������x�$��@=yЦ������w�%�$BZ��˝��B��@�.�.䫃�C��N�n���%��?�%���nnn04�Kq�>�i�*��t\�`.̟��Q�\���П��47�wi-�=��͵���ˇ�2�L��8�`�O?�8s�E+��J`�Ե�/������ς���G\j���@s3�5[��{呰��EP 7�q_t3��fc�G���3`�	��؂*�nB�$6S�]�0��R��9)I+�i�[�b�
(�g��pIE�%�`�6��j:(k"�6/�sM<�,A?oX�w���@T���7�p�x�>��C ���%��f�0+T�87�����P�� �|L���&ф��%����Kؠ�`����0g�z��L�̗�
�ܠ����#(����p�VE�E+	e�	�$�d�߷�*�h��c��0Ի��v@��)���3�b)z:W��u�zo�'G?Il=��KtV��(C�Q*�'���PӅ&���s;�� �b���7�~������n���9���s���-��g�r�Yj��)*��A���y�n�06ݧ^�.�X�m���'��,r��S�:8όR'��Y��$46� T�"�����@˨
�kg�B<u+����M�6�Y�0XN�����J�Je��:�D�k1E�𝺑:Am�Gp�b�ڿS���q�7�.����ׅ�*�0�4|�5x־��(��d���n��C��3��P���X�	��'@��zE��;������aͿ������6�*]H7��77���C�2���S 7��q��Z��2�/uh��ض��&ԗ��AO�!�v��_A��������R(�����
�jp��!�B�>]�׃6��/3��	�P�*��o��q�t,�z>A[�^ O=+������5�%P�4�+��A�A�z����^��!Ȯ���q��k��p����_���å?!�߉�{�74�K������'�4�p)
����h�� ѻ
n�"�2��L�V!0-g�iJfG�ٶ� e7�=3�a�7�`|`N�������9��c�\ZX�i�4�J'��!H�i:M�$t�9`5�⢄Ϩ!1�fa���QL;��� 4s��;Rp5���{�T(����<���2Z#�(-*#�v�N�^\�%�y���&��_�P�kl�>�1���ݏ�	+/&��ݔS��K��ك�ۅ�� �y����sB�E#s���.�P��P�J87�ք3p�:�v@~��M�y8ˤ��sӠ�`?���p*�ܮ��َJC~8`�G� �4C�+r{����ȣ枠�~���������e�;�/w�����=�D��
��3���l�n�3h`�3�8�f�~]Ce��i����Rȣ�7�EX4�U��+I|Dԥ�F-��M2ԇ��{,$�8>�;<���7�X��TE6�E�l݊o���=L>�eQ��>ST�9�E&�_Ē��d�}O(��W��s���|�U�=M�򰞉���ZQw�{���IH���:������Kk�R�qy�_�\����׺�����:b���F�=w��ү�NK��������1���T�7px�.('K���������_����߃�L�R�r�����7�+�9Ͽϻ0��R�y6�E�S�?/��;-����q�@�A\�!O[!Om����/�����g�����Q��`1��">ڊH@4�)���o?�M͝+�|�	5��(S�=:/�S��Fܘ�uMDQ�i���"&_�jg�{e!.�oLPOb%�N?� b�~���ugwB���͜7����ӂtV����o:�8dy���C��f�3:W���y�P�#,���w�~O���]��}���gق�������?�K�O������{�P�}������&0������[�M�l��ˉ�U4wكٿ���[htR�s��4{�G=��I��@Od�j}�z�x	��9�}g�k"j3�~G���Օ��s*/,:�e���x����Z.���:�Pp:��Q&�nv��a%��R؃c3�����S�b�g�r��������Ta�0�1������<�K�8���r`l1L$�
�Fz#�k�ݏ��Lc
0�1x�6L��ˉ}�-Ʈ��c���aF�c=�F��n�6���P�0�(Vˈ��hb��kA^�����a/c�0��c�fl
V; ��c�R�����&���Za�b�b{��!��WX���t�!���0D�5�G�6�Fj�g��pβ�3�>ȿKÚ�^��D�
ZD4�B��h��KA����~�m�*�4�Z����ȄR ���EO��Gc&�l��;���Pv=�*JX�*�Pzm�B��8 �P"�y��#r�zoi��gNpC�L�����'R�����ιeh#���`o?Ț@f��$"`y�����u��1�!@�	���X���}
�e/*��m {����Y�q�9L���@��D�_г���rH[8hᄛ�'Ч�	��{�A�Ehs8�;m���(w@Wd�Z��CB��|?����F Qk>#�k>w� E �Bڑ[;b�D#d���4�K`��F�{�����|�"m��Z��i�Y���;��-Ї�"�Q:�H֬}K(��ǵ(��
��gu���Y�D���'�́�����?��E�蟢{)��sլ&���i���������
��/z��q�Aܵ��w�F�V��;��ڟ�}u0���$ү}��1�g�'�%G�>xM����J�L�=䎋����5�
�F��g�NY$�ܝռ�_��Z|���o������ǽ]�omI�T���ӛ��=�7���qe5�MS���uc�V~a�"[<��C*�9f֖�Ϯ��w��:}o�p�J�o��9���Cή^J>�=w6�QmxN�XTO3�;Hu�c?I*a~��~˒.�.����'/-ս�;�v�����NU�=��e��b02�w~m5,x�v�ei�!/%�4{�Z�qv��8�����^\�"�̹&�����\C�3����]9&�y(^+ ,�����kodG=>^�Uf/U4=6vBUM�,cS$��ݝb?�W�"�=*r�0���X��k��	(+��c�x�Zd�<^s�����	�V����;Ƽv�
��k\2ޗ�����O�w�y�$U���җ�^��YԨ���-���nR�R���E��~����"v����>��SI��Z��%�l�1����ۇ��B�3V��G���Թ��˷Vc�O�N��y��圊_�r��v�!�p��L��e�Z}�����,+{� ���qM�+�ظ�2o=�u��Ų@l��!�y�f�E�z2��uF�p���zK27c]���&�q�"?�����BG����8t���'��z�c	f�g����1�]I�\����M�&�Q�gTR�Vk��=޶T���������+R�:Um����N���2�r4'�#>�4���r�&6�8�\P_���*���,_���g�_��x��	���;��W�h�jŨ!�N�������&-�q0�q,>����hn*�ψ��#��Ǽ7�z��D����m�ؗ�����X9�z?u>���S��� Fr(Qh�6�f�vJ!d�Z���Ɣ��4���-1�V�9:S�Kt.1����͏�S6U�y�W�E*�k�����9��*��EWM��Ǽ����s�k�i���mw�Qw��+,�~�Vo�xP�d����\��M�#�α�v��CxQ��˚��m��!uF�!N�Eϣ���yZ��L�1-��ƚrL���T꼆I�#�`�n[sU�M�Ggl)�vW�"�Ӓ���T��'B��z7����^�����[��Ǔ�j��a�P�d�Z~)L�x��q������	������e����D�Y}��*"a��*��}�_��)D��tL�v�*��*��e��ʌ�3�l;���n���oJgӊQ�㋙�/��l3�� ]Q ^�P�x��s�
�J��~'S
�'4[80���xTnRfϡN��9���x�qO+��{o�Yژ�e5>-�qp�io������ۃڑ{su�Vr��NJ�=�|��v�4c0�����;�����e�1$��љ!k�F5F��	c{�[m��k>��]��H�=��l��ކ_S�l�0Y�O��m�����&=�KgbsD'o^�p�{C��xw\�?B^�FUڗ�^��x��q�w鮜��O�U�+/�[�S�?9����A�fS�;��׎��>�(���~	u
�*?�"���ry[�2�J���/�%�9��6^����Un��2�)����v������>�0����V��Up�a?�n�¤� ^nFo��S-����\�O���ti'/*�'D�<�f�������cVϽ��c��of~Ĳ���#��^�&3eWJh�u^l�x�X�\�ivd�?���L\�q!��n\��o�Q�����R���o7�?I����M�$����j����q����Ñ���j�	����Ȏ#G��2�(���V�	��Dq����T.���C�y�x�%��O�x���Q
��~Ѓ����6u�7}����Xdgs]s2��q5�wA�.C��G��;���a&<vJ�j;��?9��9m�{0��rh��X��;��i�ۛpD.�C	6�{|� ϡ�3��'h|��\�1��Lsl�֥�q��h,�jo�6]r��N��UA���(�g'���#�o.	^����ukTI�>��)4�,)��N-��I��Ǫ1z��:M�~@ R��:<m��bjo�\�,����7)vм��*\ŭ�Ϟ�����|<9��N�oٮ�Kگ�NQ�;�2�i.>>γ�[��ku� s���5+ū&*��=5�+(N�3������8�</��Miy.,���$��{3�)��?��n4Ұ��i�U�p�fos��s����N��\f�W�mW6U��tf>uU�Q7����Hx��l2��A��e�=���O�Y<�8�Z�Y�pNG�|��9ل���Y�����7���6c?�=���R^~Z���F��+���Z/.�n�c�5�lݦϷ���'��M��"�r��*�?s��O�`g��)T����cw~����c�ă��P�9�B�Q�X�,�<���W�Ē�#;��L��(��^�y�B�ab}�U\�g��њ|�t�fQ���_H�*��?��}�ň�Ç�4\�k,�;�RO��?��u�{���a{��)J�R��	c����2�>��ڂ{w�����
�oBU�����*�YR�1���z�M0�r����UŽ��{���I�Z`�Y�v�R��D�.��/��H	���8�H��̉��򟈓
��+q��z�|�.�{�4F�����������u���u-0
[>�)S��ZO�F��}�����x�n���q>=�!��gK�J�.igAg_7>�nk�_@�&��6#����d�ǫ��Ѝ?*'>���pަ�s��Ϊ���#���,�s���a�W�E�,��9K�9X���|��W�K��[`�~lU����ks{/=�Jj����őL�$B�	�`�`�H�`�e?�]���\C���+�{�e�n� �χx����䘽��tF��j��NV�=ֳe�����sW64����_cՄ3۶w���c��f��w8I�ս�]>�ǟ��7�p/�k=�\�ب�	�z��m�;d�DdGW�W��l�]9j�(����Z���oIk�eh3㕚םn�{��20���j4�mJ9؊����h�Z=�������o�ɱ:G��eﶲ�1�y��<gA#����9N��m#"���vǖf��s�J�vM��=���o����7�%���ҹ�qԮ�gZc�ӳ�nT���Zd�DVVm�u(�p,���
�Z�A�xa�ԛ)u��奩L���W����Ǎ�`��#?�?�~t�E�G[NiG^o[7#R�ݙ+�Y*���F�8�k؄㏭e���t!���Ƚi�d����������i����,��j����c�H�8��t =������oiu�3�������aC�s1��kT�����.G��"����Α0J9=+���s����d*i4%?����.������z�3��5�|��!_�Z���i
!�q��aA����vço۬����M�gStR�y�c͡�v�F����f�U�e�"���8����W]b`��2�f��(4�v���H\�9�� c_�sE����.\�m6|D^�ͮ��=���D.j���qE�I����}\�ʱې����@m$ґ߽�����u��xF}w�����H���Ɯ�y��d�BEV�<N�1�8�ꂈ6M�3��YF����v���,�Sp�'H�Eq�Dգ���4��;T�����ҿ�z��!^+�l@��S�7�8WW�y�4��g���յ�K[O�����S���>Ft~{D�[x˨�Yz?{q'Ɂ��z(��ox�\�g׎�;'hk
�کc�q�eP�%̦?���R���s��[�Nbz�w�"�v~S8�p���C��Zx�^��>n�Z��R%���^�m_W����~�� �k���V�;�@���#6B<��I�My�#F���zY�9i,>�]1�9֨i��*���Czݺ���w�	������I~LVS�±Z�ݖ���<r;'|l�Iά#uo:Gr[SG��mV�	aK�6Vi{xŖ}���^�ض�����P�h8�잫Bޮ�����N�L��\�>x������)N�yI1\�1�}�b��4����Ş�ږ��=�u������!Ï*�W�-�c�3��s���jP�k�}�u���и��ugs�o�g����6ov>F������^n��6��쵻K�̦���Ayp��z�G�^�Ӛ�|�-�j;bv,��zg�v���5����w;'��	Rj��r\y*��¹�N5{�n.����>��_���x4����\8�ӿ��ǉs�"��$��UWR}ܨ�@T�Z���C�l}E��3=؍*���Ϲy{r7UK�Y�'Qak�C�h9lG���.�z���청ΈL:�����KQ�!aނ�矹6��ao�"5u��OW�����x��2��r`鑔�7{��x|�K�"N�ڭS$G�m|�	R˸-��~ٍ�؍jv+���q>7"�����_~9x�~��\��y�k/��F��
��1�/�������G�G�Nh+�Ԏȟއ�#?D�ԵQ���~���Pj�tsD<�{֐���/��Q�>�j�&[�j��?58��d���nq��Ô`3Zݶ\gR����x��fYk��̬�.�JR�;I�cj�F���UIA�o�;tΗ\�יm��T_�j��ˣ����rz.}�[�uu17~O����o!�!��M��a�3��7O�c%����]|s���E-�O�_N4m.�b�w�v'�pL�5W,%�,Iο�q�r��7���;��D+XM��gF��0z�iiv�T�'�����|+p=*aF)?�q[D��Jd O+�l5�լ��T��������1�L�y���N���9�^�13N�*�SSg�9������+��޺ұ��w6	���O�Pƽ�����84�o?V�E����_�~�/�E����_�~�/�E����_�~�/�E������D�C��Es39�����Q����p�7����/ ���,��	��ސM�/`f�~�W�����i�����NWI��/%U�$������a'��3�筤��Y�w�o���޿������>MI:/�w�Oe�K�$�����ge�L����[�s������o������dȩǀF2 ��ô��K�c*�1N�Y���f�[8�se��WkU��~��@/�		���Ȕ�Kr
��<j�~�! �C�aK�f�)�w��eYO�[?��t|��T�E��-��#3��s}��3p18�Ԛ���E�59�4:��A�,h*$;$/~hwp����Uڀ� ��zJ�׈֖V��`[�u�x�	�Z�!��={�� zΓ��)�Z�,(d����C,깬%���� �v�� [�;|A��Qa���dk���h������������Xxr�ɬ��<���y�E���NA�k͡��c��,Rdm eJ�媆2ȈX?�ת�!<P���~*L�mk{Va�d�:���a���tiE~��Z�k��D�P�����W=�&P͗���� z8�Š#�, Kz�,剴d���W�a���Q�9=�UOz�^�Om��YW<��p�Bo�WN��������.{�����BۺC����f�q	϶5۝�<ȡ�5�]z�9?���ZC�a�v�s=mM�A����
m��D1Sԡ���ܒ�>����z��n����m�h������K����p��6�����0s>�jn�xK�*_�X��7�0�VoMf�J���JRd����B[-�X�[�A[agi�͵U���"��Eo�0�0��,�z����E����O��gz/0�e�¸�G�)�4�U��9��Ō���}*�n���l����@~��e=��U�Eok��E�r���b�����2�.���9E0�������az�2s��}�Z��j`s�v����t�r)�_Ơ:;�4�/�z�A����@����J���~̞���N��L����:@�U$��-p��������@�Ṷr��Gr~\� ����?H󧔦�o)MMg �r�������s�ͥ�~��I�I��8��!/%�54f㚚����`{V[s����fzjN܌��B-��󉤹Dҟ'f۪1K`���lt���4u������Y�k�B����;�W��`}ޱCZBz�߆�� �n`�/��H#�w?/�񙾺��y�-��wRC>�w ug�1;�x����sr��-��k���K�۫�#s�z�9�ė̗���2����>��/3���>�W�2 �����%���{6͇lEso8^<�����-3�.�k>��:�o�n(B������]zs=���;��ma��8�ʟ������;ɇ|~�Nr:��]�3-���Ut#��[͔"+�&J���
�
����_p_���o{1.bŽE�`X �]B���w��Uf����0Y��A80�r<�������	=���)�bA"9�[���I6�v���+���z�U�f��ӵU^l���ȸ4�"+RWO����;�b��9,�����9[�fs{<KcK�6����D��j���G�+��L�����SX�2T���	��O#���w'���([�0-uw�Fݪ�7G�lS^�9���f6�T���B\�X<Ji��a�X*�j��!���[#qJ�3k6��"�)�-=A��{���=�8��w�R�5�)�C:wk��v%��gL�'�ٟ?,~9�V������l5�z��k��`:��B�MTs�Kn5E3_-�8�aT�aBS�p3��{��ǋ��2b],�^�������� �dVVn��/~"o��aj]����J�%���3ꫜ���g]����f�gt��e�9��.tz+��bU���1���.v�;�?竵�띨+��[y��b�9�>�m�Ci�Z�l��;�$�K*_���]zW(����Λ�Դo?���*���M;2ۦ���s�����/���z�T\d��P��};�U�d#��i;χ�e�H.��X�ͪ�!��j_#o��H�����괩���n�K������Ҵ{�g�bظ����X�w�=��ͳ�xc�2�(|���n�7v���Z՜���J���n*^^Y��J�־l��Pu��j��ᕾdt�~T������N���r�a�*�7�$x=�o⿚�S�U��\(�p)��`a��h�l֋�ra�2�咮ؓ{��
QΆqi�
�r��O#b<����Bo���^Z~�Xo�FL ��R]I�킒,��M��<�74�B����%���=/�mb�s�5醶�S���>I���{�Vx�.TNvGxo�M7��4Oy���e��S+�#��f�D��wi>��Į"D�����M�;�N�l{�wu�P�㨦Mo�g����􎈉�3l����_�䡲/���+�N����N>���[M�0����Ҫs7�5�tS��W2�k�
�iZ]Y�y��W)�\f���أ�Z��Z��I�8��v��e�m��z|���O���#�7�MZUǵ�?:LfX�T`lu^��U6��ɠ��;p�"���N���a����@��l�h�ع�����/-��&��Z6�dwF<�r<R�g�&ֶ�f/���;�'��Y�����,~���eieo�E{�S몫W�E�q]V��629�g��#6Qk�Ja�����i�/K�$(�����4ާ8�|���cR��o�gN<��y��={�Q���&�Il<��o�v��������ex0�� ��S�z�;/�2Y�-�����h���p�B[vf:��s��37^��j~蟶sp4vdu�a݁�7W�BN]����F�8MY?��L�G��s�hyU��~��~���Y1��X��RN�n����^�|�C����Z
�E
>Y��l?拪��WX�}�6R���(���TS����6����O��go�T�>��
�Z�
�_����	��в_��¯��M@�_ާ-I��b��n�b��kW�e��i�vY�&<�F��RZ�|����zIhj��9ԕ����%=49M�2ٳ1��7���j���Q��a��vro�nQ�n�����H�;��	�E:Jd�븝;�o(�<N2~; ���q�)���0��Ѧv��;�w�&/��o3�}vj�큔��Ϻ����ϴ�^SX�f�]ۖ�y����7��<��;����k��\o�:�<c���&�OJ���~���0%�xM�k���ٯ�p㴫�!���t��4���KR>�56~�QSzU��5QE�79{�vq} �s���
s˼��=z	2}9��/Y�I�tt����{^�ĩ�ݷ����#�F��{Sf6�µᅔ1��l��:-�ÎG�M�|���$�n��w��{3�%Q�4[	���rG�!��zB]A�M�T��)��ȴ=��e�y�zx�ɪ�e\�����_�w�g���C������LWyo�T�_��f���!�+�$}�G��=�X���U�oN��&3���	��[Bw�ěV��.i�����٭t����լ|����qǎ-fX.�M�|2����ˡWu�E�;�W�����?�Р�!L�+�^^o�^Uw@��֙��RW�u䙰�ɑ]��[��ps��򀰡f�m���}VqJ�T�����L9`�j3�������9;��v��"or���7��}�ݶ�S��]�����t�k)��t�x-c��J�٫3_��0؜?�&O@
��3���X'�z��-�������O#O_|s�yݖKg��P�
4�p��d2Kda�foݫ�������y*�!է��_Pz;��wĿb%?Q*9=B3b����N½ʍ��\c��N\u�a�����\���V�:�`&K97>���z�Ek��a��C7O-]\y��u�D�D�èR�1�f�w�<���KKz����U� �ݡg�w��DeG����)�-$�qua�B�{�.9Ӵ�Z��j�{���U�ܗ/̽��\MߍuWr�%m�o�د�����cE�7"�w��7��)߿��'N��D���܆�٘�*s���g'O���Υt�̒����npQzgH߉n±�I�Ux���n�'ܶ�=zI��`��4��9�c��,��:M�}���u^�N�m:^Wm���n=���Z�{P�I�^ ��s���"����*}���)��
'�������rȚg�.�@�;����.�8�z�ٍI��9�О��W#=ǵ㟻�o��_:e7V/*�8��O����x]"��2i�D�G�y�WQ���Q�R�]�/7?�i�V����m� �N���u�o�y��D4�j�N�w����7��C�Ɩ�4qج5{�,��fV�k��$5�E���+��ܯ�t�����d�Ա�W�����Wq��������d.v�+yG%��n~��;b���d���'�ų����o(�����#EԀ�c�
�'��ʧ�N5���/��'��;���g�����Ӆ���¯*=�jqu{���z/�1�~��`nߢ7��O=�LH1P����t�2�*�c"֞L����mك�K��q�5��I�x��ո�ш��z��&V|���L<y'{����]�M^��ݑ�^C�dH�UE�p������{��q��rđ﫲�z�˿��^b7���lݜqKS�Ϟ�.U�7���J{~��� �W|Cy�d�Cw������!q�Bm:�1��}��<c[���,|i��ɭ����}�cn��)��}M8 ���~�^��`�^�0v��i5z�>O�;K���'qO��E�$�/�>�-#.3��{D4���y������5�Q�D�3�/�OaG�C��;��1]V���:�B��/?�_��\὾p¯�Ɣ^ԛ婃�CV�jE~U��.�~O*�(�b�y�|h�3�KL��>m[���������~甎o��j�ZcZ*"�0�$�a�c�8&�+�����#��y�pc���=�%����ݘkh�b�%���o��z}���?3���<��ఘ^��d��j�5�������c�E=.�g���q���Ҩ̋��;��G�[��/�����ې%��31���+�m(x�'�K�A��o�4i��3~��kJ�X��߅p�OQ�C;���_NP������?�*�L�h��4�`CD|�ڧ&F]�$>���J5p|5�]H8�}��dOw�f��Wwo�����NC^l��-Kn_����p�y@VH���0g�N��뮚v��Z��K���CpF<��|�⚿����
t,�kҾY���p9���U����B���x�!�:~�#mo��F����K��`�o��{�y��1���eRi�y��y�W�{�>�l��L�/���������m�]3��@�Ⱦ���E�u�ϥ9=��exce�����W�� ֚3{>f9J/y}A�R܀�=�B��Ÿ喝���B���_^���RZ ����ǹ�>gr*��Y{�s1"tob�}QU��Κ�C��_H��nm���R��e��3��5n�*�TGD���/4w[�2�np�~�/������̥���V{���C���"I=X&Q�(�m�����ʪ 9���.�F+���o]�5Zn,������������b��8����*&�e�͈��OͻW_]�9�]}��J�CqRvn�˓�p<�US{������>���N4m�A�^��ia�z	˿Y7����PQ\'�u�n]V9��Tzv�n�<�[ߗl�-��&nd�h�vQ}�j��O�oD�t&,�`9�Z���]LB�"O��m�Zf�+S�6[��d������3R�E���*�]��=�{K�yA���KW��*M'�Zk��YNq�I�>j��p����w4{S���ANwoю�i6<�!:l�J�U�f�n����rⰄRd�3����컏��T�豈^����P���ǀ-@�w%S��2Q�%�sLP���G�I^R���r-VMf�%�V�بCW�:y�����o�LW������Ke�Y���n�|ɖZ�[-3�c��@�t��Z�sɇ7ղ�5���|���W���z'������x5��٢�'���.�e�?�rQOh�ճ�>�}yKn��:X({KI8:~��gH�+�!�&Q}������d���q�Q��5*�+o5=0
}��V�t����D��
'���Q�Q:�[��[��n�	�*0��d2����l���b��[Å��/)�_����^4+�;������Q���l¿rs���b�	7�K,�����5�.����&��^�^��59��
+_]Q�<G��\;�㕳'�ѹ��9��-��x����|�ژU����ǂ�vlV��g�q�S��yȋ����}�����{^E�2^;}v�"N^�}lO3�B"���Q�L��Br2Zn�x�z��c�r���x�紕�ؾ�:��58#�$�2�x�e���Y<��]�벻�:!�}_]!烰��`�k��_|T�S_߸��I��6���Zm�F嘆<�>
''z��/kE����O(��2عo���}k�^����4�R;�i���V�ƝS�{�Y>�z��U~�ɍƊm9*��&��
.�����"^��v�g�a��D����S�"'GOwu�8�3L	�e��N�6UK���P�t$p��ت��&��ݮ�$�c��ԁg��kE���f4X ���à�C����Npwwww�ww���.���$������^^UWuU_��e���6���L�$��]�	�F5N�4Q�ꄛ:�BH�؞-V�@�#IزVyKnψ��@�WmL�F��ș$�����cлG��c����ӲS��������=��Ǉ����&�+���r
bz1��D.s[K�~�Ṥ���q�t�{��=(�m6��M�@>K�MhG�Q�r�!c�#�DUL����3�kMG9;Xj�G�$k�NՁ�)�P�|��'+V�ն�iU�ߟ�n�8R\jE�9<V;�?R\��WU[=v�L��Q}����.�HG��oʅ�=�ȟZ?:\2�
ly��!J(B���IIH:�M�dXV���]����.�\�2]�gm)<Y����X���6�gm��L_�}� �R�Ų�`6�C����#an�ӓ6tuw^�a�3�5�|������~�vF.x���������'P#�ȬW�|�[����A�|��-�9�����g���U�3o�0�i��O3~Dw��#����$:U+�Ls�X�R)�^���(>�%��v��)�[_�`S�@�)|�;d��V�{h�������S��^�y��b�*�K>z��"}�!܄]�m�UÕ��G����}�
	�6qR�>����I�z�i��-!֒Rh���,�'����R �5�L5��HjG^=��X:��	�y�X����ʆ�{��� �-q^kћɍ�Y1��&��g^����gf˪��=��y{��_�|c����)�+����ڷ��6�)WR�R�X��>,�������?qWi1��f������;':�v�B���\w0j᜿��:����mHW�N4| ��ņ#��HÞbg^A�.��gq� ZWW�Z��KGgGeF�^m�GDx\�І���H�r� ;^����3��:��N��#G�d[jU�
#��,����B�Px����f�a���bk��q~b�%�*q�iV7��Z��p����I�0f���JMTT3���x��\pPQ��a�wj������LLL�]��WWx��~,֒h:���Z)��9����	]�ưy��@�Q�m'?�@�u��7��|=�G���$C�f#�d�l�V��w��� ��q&� /����ƨ@LM~�4�O`d��v!s�7!�!�2&�yV����f��Z�YH�F��L~��ξ/�T��G|RI�ejVȱ���;>���6hbqi���W��n.R�,`�c5�;���.����kg\#-�K0k��	�K�-���7��^�[����߉2�<�6��$�XE������0ʫe�T�������P-������X�[�1�6$�g�%^
W�MWO*��Aу1%�1���Z�q( ��m�	Z���3�^#��(duU&d�$ѨF*l�[�ID`�K��(y6��H�I	x	㶖3���� O(���+HD
�]��;��b�	��S. ���8�[�M?��'�<�;lF[sR-�p�l_�@I��j���V�N\���KThKj��o�߅���&:x�0�nM�W%��蘔��*
Y�~�\q�j]�0�Y6C�,G���=�;����c0�C�ʾ���G��K��B�x�Ӌ��e�S�Jp�3_��cg8A��z�eD����0��w��>�_�V��
% G�=b2���9��q�*��H&�Ӯ����pg��ܙ�e���G���Ԝ��ʚ�U�'�mK?
��y�����;�U�T��x���/%�i}�V� �y0��Fq���^F�.7�zK�EbI�rH�>V70�E~��HyL������:�7$���=%b��k!�i	��]aG_%�ٓ���]��9.�����x��`�p�\�}l=�� �-3I��3[M��I0n���*[�z{ִ!�^��[%����@���j�q��&���=�L�
rO�M3�f6VE��!��L�@�ȱ����֙K��v��ӹ�����;���H��j-_�.��p��:����"1'���<>kn�C+���[,����KO�K�Ί��AG=�+>9��d�T��.���"9�%�^�6�,H�o��:�8�9��a���1�77��*b��Zi�k|��%f�t�VT��doQ(��`���X|Gɑ��<$�1�*/%�*b�J}&��u�X��z��/� 3?]��=m�H������b�{��)���^8�#��Kx�Rú�WZ�F�deA})�_˓q�P����#�߹�(���������e�{��'���XJ<"��a%�Ѩ���|��f�[��cT��-�R�a�U�fLX_��*V�C����3SlF�w�v]I����_kr�N��$7�p�!�b���H�U��I����)��04���i��@��)&��deа�'U(01e�67ch�yM��*-�:qz2�1@;�&k�oɪ��H�A+����0�*�(��P|�Y>���ny������6��p��:Nt�#n~�UOG�	 �lůϼGb|��A;��h�T��Y��Í�bD��ηsh�:�ጣ���_�|C�Tww��ZdwSҺnmb͛'��6v��߱*��ٌ�&Av��K�ɸ*�/l��-��������$rT��v�J�;x��&=V�n�`��D{Ͱ�j��=��������}'���y*T��[�_&�?�S��j)LB���G^u�i+?�i#g�e�Υ�ΏNd�Տ5�6�Ԃ��t�k�����}�Rv�����l�IʹAö�z�u�����J�'#�g�f��.n��*(E�����}�g��(>�&ݶ���}����CNpˤX�M�B$��PFi�G�f��,�Kt449�V��a��w���k�S\� 2�1�s��y`Jl`�9��3V�#�6�[�nn-~��4��a���-�B�p \��XUO��:�)��%rv��#$��Ջ_W=)#n3x칚���?��uVGn��[N��7�X�G��_W�����7����V�w�`��-�Q�J���jJ!� �2���6���\� ��A�x�\��r���*�K"��i
��cg����%*�^�"[%���e)�_�	K��/�a̗�7A\�a�`,T��)W`*]ʧ��m�J���ש�Q��*��5�-</��
�v<�D^t��J�_r��[��t��Us�K���ޝP2nS�i�2�y{u;�7&Wu��0�ŔE,�L�C.�/�D(t��	j�X{J�l8�|T4|ְ6��.6�=U铲X��au�l;���_}�G�ۨ_�E�K�q�%j�:uGi�2_6o�+�F2��?�֋+mW��B|�Cj��{2�F��K�3v��zY&�1a�_�Fzx�I}��nu��/>R�ҳhȢ���T����� ��3�N+÷ڎp����DX�
�����(�D�ƺ���G�"��\�iH3:z��^�Skde$�>�A��͖L���}�z����(�l�]��8c�E��
g�����K�6�t4n�l���5N��Ĳtߣ`�%-4�X���-�Y�jsw������Ñtض½ȖH6�9e�Vʭv4:��ޞ7��n;"��(�+�Ⱥ�Gӆ2��L��"���nW[vBŭ���u� <	ԚjE<�����������G�7p"���l�U����IM�(�\���h��B��x�0�O�Y��
����c��#�6��~���qV��k�,el�\dx��V4
�q}) �F��V��f	�{�������:���Y����צ�0OS�TS#E��������6{��jZ�- G�[���Z75!�R��[f8?3�-����%Hy`����DBy�֏k��܉�'Z�nf�ȔD��v�f��τ�y#��\F�I�N���u��0���u�St�MYl�\~�Nl԰TI�ܳX����h
g��>�L��������,o͜`	��%���$5ŷrUa���Z81�9�j���a�B�pM����:�e�u�9����UIђ��2m?t�`�����Hvx���}�_I4���y��mw������y���fz��V<v8�fvmiX�8k�V��k��x1eRz r(�U��[���9�j�����R?P�\��y�Y#�����K=*��h�5�'u�-���7M�l0N�u��"���-��#�*e4g�%��L,|v�V�� C9�M�v�d��\��Q�+,�j64��%�F�L�^M�M�ۻ�vz|���n�3Y�9_c�(�Z���K%gԭ7a����s�6�Ś3Y>7߷�6�l������x0#�6�,�)���(~�L[]�'�w^*���*��+@f9�>��K��������b��0�[����d�=���O_U[+���>#u�����"}�*�s{�J�W��"����\�YZ��d�ŀ(�B4a?��O]�����F8�P�O��0��P}2
��ԸI�	���F������7��΅�է�(�¦���>E���h��+��結��GgkS2K�]YeF���i��=���%|�j�3V{|Ǒ��պʯEx.q��7w:��]ؽ\$���mҖ�Fs���ڊc��Ys-���Nm&��n>�_�}�k�;������!![�d\��%)X���W&���y[��k���zf��ٜ�\(�a ��~X�.W�{]F=�;"i�Lh��D���]��J+w�&�s˔9� �-�	��j!�9Ȇ]���AG�\)_�W��9,j����.(63�떇�a���#e���)f/��ȴD8�=��	I͞�ݧ[ϭ7r�y�2.�1�>��#0��Ю��d����yS}��}�Yh���F��ͧ���b[䚯��f��p�ˈ"��֍��W�L2A^��g�H�b����մd�qJ!Ҝ��;���<Ӊ@קxF� �j?ݬ��]�4_tgi8�m���Q��R�rcg ��A��;k7}��;��"�E�V� b�u.6<i�y���[E��
��!K��+<�;g=�^S=o��Iv���v&� Ʈo���v�~cP���rѓQ)��4)�i|`�}��MR�ܿ\��B2�30t	7z������xA�2��!^�1U�V�?1�D�Q��"G����cr�[ ���Yp�7�ϻ�����Neo����_8�<61��}lli��#�y�~��V�J����dڭ�du�uM5!,�IEB!��5@�Wb�\?���tE�0��!A"�F�&�hrYn ����	iĝ�)���`�pzl�K�\վ?�%cOds�ڲVs�p-8�D,�ڝd<����y�
�_�H�9�z�T>�ߤ���y���߇� �85�O�#�}�	pS��VA�L������]�q��8��L�Lh�(�cE�C�2��`$`y��iM�����}'�Re�NP$jfj�Ri��������J$眱'ZƓ�"ρ�\>���v�Φ`i�b���ܫB����t�gӍ�*��6��T#�0�E`�a�Ⓢ&�=��t�e�wm�#�?NS��+���Y&6X�M%��)"
��<�M�DD*~��/��u��V�V���tX�M�������:��'�I6�{$u�TG��#�:��T$%��.�5%I��W9��pVk��I�`'_�A�Y�6���y$���(0oT���}� �3�1����K�d���=�}��`z���o���C�z��,�ץ��wQ��`�=k�"?	4��J�=�h��]u)��O�z�@Ů։��3<��Q`�ᘔ�%ıt"�<ZD|���~���XMQ)˙I	&P���Z�����YehxTs��p�+�R(�x�x70��F�B}'�����Ehz&�48Lkd{��}�K��+����3���J
D.2�=�>����E1�o��I��90�W����"��i��P�.7C��'�!���a�Y���+��r:�۶U���>����),"�G��PFG|�n�0��u�:
�ܒ���L�6.CR��U�Γ�+1&�F��@������{3��><E'�k����c�z5��Kcx"���Ƣ>X��z��ژ]V@�6�g��)W����D��ut-�|�����y���m��= ͐�9mF�o��P��a��;�~�L�Q��py(�;�G�H[z�^b~��>�)'U�4����`����)<�^f��W��Dx���CmH���ܣ��Iw�Vd�hF�	�oAʨ8$��`p(�����VIb�W
�N�4�Y}�������/�g]J�v���p�QU1+I�}a��p�|�J<�#&*�5zZBy}���������zn��H0����n�qFq�k�TM.YכS԰ֻSx�,K��V�ג��謇�ka�0]G��^t�P���-�R���Q����Qj��o�,8lA���Ҩ�%�N�y���h��Ú�XE��]���Zݟ��z�SJj�k <�f��a��Ԯ �MD�O�O����9�N�7���=��3�U&Ql��m�w�TBC�B�T>��T0U�C%��׉��|�)�ۏ=wZ��P�v���v�з��̓�^��+�d*x�������c0�0�����`��>��O���������G��O�M@�MDL�BM������+����o��UX�.�\�������Z9�i/��'��c�jAi��9_<3�D��#���*qP��'t0�b��h�t�9|Oj�^s~�U*?�oQ�pmO�74E�s�"`�Y,�~("j�`��ވoײ?���t;��QZ�/���~޶3s�\{,s=�
�k�q�v$Œ���PrH��SP��i����H�o4��Ā�Jx�~��F*��!��j���P�����P�2�Ե���$�;b�'��H�o���mW�<���L^ז��RZd��S*I
Hl�����ܿ%�
X�&�&>L9�����G�S]�f��<�Ǐ���!n*�t�d����"�o�4Q��x��7����lo$P�T�U�ҟ�-�!�m�901����\�������Xo�[��y�R�b��y��Tbʟ��{��<#\���=`�	�Y�8e�t��Lx0͒���,B��I�g۸����l�ԐL�\�"�md�'�Yw�v�	9�M���r�(a�%�����7��7sm��݈��K�6߬zP�W��H���H�0a�$�e�*����|;�[ ������C֢*yzaJ
�R:Ho*Z&�s�o�2�O��f7���.g�B<~n>�#�r懐��U^,d+����IȎ�
yh�x9K�kv�����܃������0�f������0�0A������j���ǴIU{�=��-��L :�.F���u�[�N�3S�l��y�����Ɗ��I�^-��^�����ԇ���1#�f:�\�D}��Ȑ���_}����E��]���&�1߫�>�<�v�9�d�B#�v�L�kό��q&0�4z}�����ET&���l$�ٲ���?"��aûB�~}�7���z@��p�ĥަ��Ci*�?Fw�dx�즹������C��m�Z��������v�����_8��t�����+=5Ȝ��?j���m?��s�?^�W�s�qb ��>�k�g� ���Up)߽�Z��?$����z?���
��3t���Y�R��)����4GUb$��i�IrQ�&>��	J�Q����҆�Ίl��|��/9�6��f@c�v2rS���)zg�:���~���?t�r��}e�I���4��/t~j�黯���l�_����-�n���X܇)�S*o� Rʺ�3)��������΃z1�f��W^����.�}�&��X �$	h@���RW5�唚�F9D�&e��l�!��z����w.�Nh0c�ȗ�NnZ�bK��L�j��f"��M{:�J՟ȗ���Y��;~��
�A(�ֹ�&ۼ����
�13/�9�ֽ�;�8mK��6|�$�x���L�A*���1�eE��b�Wֽ��>1��p|D�&��F��Bs������A>�N&�N|�Z�,\�(��<Sk�
H�vLj�>�J�����:���c�yW��~^�����0ᔍ��������_~�����j�<4���3!B�RI1����G^	�!#���<�N�"Sg �B0��B����M�%�X&`Zrd�Nz88�Мr��˺z;ȪJ�57�A>�T�wp/e�����G���W�i㣟f�K���R���8E����n�$	ҕ^�@�ml:4h��[��1�.��x{t��4fk�JZ9�|����:{�j�����_��%O��"LȀ}��e})j(��N�\�Ԝ�G��YV�El����s�p��R��1O]����5�l_�s
��MRʔ���:e����w"z�R�ӿi�`�o{����oVv�w]F�����J��y�}~'�&�R����~�w�8e�r6%�����q�O�>2�7�R}1��'�L������}wÿKCT��Z���h��;���P|&o����i9݁9�y���V�/�y�<PL,x����i ��G�dQg�O���7A�P����)Ja��ZJ�i�g3fvwwt�?EƜ>��"�A0��FS5vb�6���x�S� �PȺ�x D Mp�~�&�t"�o��x�Ĝ'6L�h�k��d���/�S����GP��v� �C�@�h���,z��Kp�::�[в�\���+�;�����S��+O��˙�`XN�$I;U�i=٬C</��t�,/L	Iv�sw��=���	6����'�u���v�p���u}S������~dܱ��p'i��1�Jt���k������~n�`�j�eR��Sԋ޹h�c߮8{��:ɔ*ƫ���Qr����j�oy`;���b�S�|/G-��D|��W!d��b�
*0�^ �
��,v}�ʩ��d%F?��fXn���m����T�7��@}*4��+>t����&���-�l��oBo��������4=o���h���Yaؙ0��\�����l����S�EJ�cI��G��F�}��Ӭ[�NU��
��f��zO�8���6_�D��/��YB=Tj0����&u�d�PC?�j	}�) ܙ������'���%H<��A���t
䌀&Bc<�|'� o_Q�_W�}*����q���Ӭ4)f~�(�>RwJ�灌cӓ��}��B�u7!�>^�����}����NW==E���
아�U��[�.�s��5���,����G�^�j���U��U��c��x�;�͎h�l�V�l
���xR�q��,������>N.B�1DPA�SY��_2���-`K�oԇ��ڰ8��VJ�G
X����و��I�G![$��L�!�8dtT�9��H���v�r0��WGo|@f\����?�-~o:�6BN&�Պ}v�x9�p5��"��/{��u�-�x����l�5�(}�"&��'
�Ƹ�܎��݉���yۋ�Kd~pj��":^t��t�Ÿ�r7�h�q�ߙ�<����W��k����[-��5���u�	��fK�-.�]il�{p
V0�^X����1�e�NF[�?��Ұ7P����Z��u�[UZ�~O�M���%��u�'T���3������	�[h�^�i"!_d?��ٕv
�%�m��`À'�Mk�x-J�@a�WE7AzT'в�S�8����Z��c�cә�Xg�,+���!�,U�=%���7��'ɨ���|�d��/ܺ>�;$ۜ��eM�Y>�����5!RP��� :�f]D�����\	.B�[�S��ie��zz-z�$�o���|G���<����ie@J���T �g漟|���v `u�kǞ�\����"/�����)��^�]Dl-�+�����s�3	�i�����y'� )(֡��d>FW)�}����.ܑLT��>�p�c�l�,{G��i����-�C3r��獷#SE�:��FLc�Tg�����sh+�f�U^�l�*"�Kco|I�J��@	�@�:�����ȉ<V�1y�]�O��T���;i�Pqw����/�y���I.����޻���"�|�3(��7峇c�*�Eb��ޣ*�����t8�I ���D��&I/�E�q��o4|����G��	��FT�+`�u����x���X��>���
����hj�#j4B�'n����F���k9�=w.�N#nP'�-��כ�5�6�Sx�E�i]	O/�ìU.a�^o& ����"c���l)Z��^���ߡ������x�A����vƬE�GC�R��Y�!�gG��m�J�6	��qp$��g��$�K��-Pt���L��|�R�S��Yp������ZCǟ�
,�ȭ���Z����R��)�J�	���%��F/�~��}��a�l��8�#��ϭ��ןS��L0��.7,�_fH� ��'��-�)��3�|ˇD��kF�������%wo��h��c�Tڣҍ���>�
��gj�+�#���1S�94�����8lY���%�&��MO������3t�~J����.43�iߥk�(�JN#�9��)�R�~�Ň��5)�U1�Ւ}i���9�l���x�3�}v��:NDb�l���y�9���:��N��q^����!wO�$���c���f��V)JW�hr\�T�Yv�L"Mq�������x�L��m0:�"y�=�o\[,f
���}��M����R7e��t�	K�jnL<�y��y���<��}G��xB?���D�D�X k�8y���ģ���J�T�ڟZvwg�M���G� �d�Rv:����?Ze-�@�1�Gܬ���F�QC�ӳ"��╉���Zȯ��5��ן:�~��b��:u�}!v��r�9���k�(����E�1@A��/�vs���&N[��\��*��A��?��z��U�;Q��(���dqF�w��f�%�uJL�}�7�JbD)'Ao�H	�����*�ʲ�R�|����g�8T�H\��~��x�f���
���*�2��	6Ԑ��I���J���Ev��0a<�7�E�۸Kw��7��Ͽ䵒��mq�ruI�9�^�(B�k�R?��g�{S��{����pJWy�H���8��Y�1�o�A:U�t 8��uzP��8J��.�/p]�a{%�7� �4��ڄ����zf��%Y��5W��*���vp$���hG^�'�1?*q�c��l�o-�`���{�Yn7�~�S�;?gjڭ�f8�����<����ɵ8s����C M����F������P�@Bb�]���X�I��<g�n%�����Y(�ډ�ڷ0,5�����W�X&�����H�b�̆�	���{�N���)bL������i��ԧy�%p�;�&C�̆t6hzC�~�n�lط��� �:�ޓ�k�<}�)�f��%��&ec
������)��L�ot;�u���|�����¡ݱ��Xe�~��>ɾu+�9L�y��qpB�"�����Ah�ʤu�l�j�A�t�?��(���M|���%��u����@m�j"
T���%�I2�<���H9�`0A�C��~���y��&�2ٰ1�6.�^��s�l�x=8�'xQ�]�I��aW�^G�9yX�*�=?cE�6�������7����s.\bj]<���Ϳ���GF�|id^�<ө�^W�[�
�w�<����r���M��H��Шß�d�3���/ �[��J��L_H�������a�.��\I���F�'O��㑘���,PYO��$���a�7iE�v��^ւ;��H�>�	�2����Ns2��"Kzs��@��Ԯ؎B x�Smw�^���)n�P��;>��yO\i�L�J��������)Yl�(&�O�X��/��&���C��6�0�<cIv�2��%e��y������Ng�}!pW�[[��$�u�7��W~]"�|�_ǁ��=���=���NX�ؓ�n�(�Ǣ�|�j9�sb�� �\�6���f�Tu���˛�^A� �J�³�I�,�w�?�����)���G`�/X���Y�WQ��V����ic���iS^L����3:����0�:����ĜĨ͆�����˂v�.)�|���>�@2���V�,ê`������.���������[%�lW⧾���B<Fe�ꓜ=�Ϧ7�N}��3<jU�ig��ٲ���N�ݚ�)����Fa�N�]Y�����k�3�Dc� 4�[׷���w$�P�^(�j��B��>�<j���;�ጄ�m}�2H�����h��~��"Ch�������=T�o���?^Q��A���Ĉk�p�������WjV��l�ⵏ;��)��Y	BHp��.�c�q�w�����w;�W���*���Cր���9ѝ�2��A�D��E������J����#}u遽�#"�A�{����������N[ޫ�)���]���I] Cʕ�*�a}z�
T�|�ք�!�Jn�G�f���h�S)P��������{?��Vj��C�
G��b��v�@� ב��T��fyk�=��M����՜FcI�?��F��5��Ǝ����6�����~Z����7q����O}������m�L��*�|L� ��)%����Z��X�b�c��M�����?�d�����lݬ� 4��5�J����A�nC{b����ϒ���ϡ^�_�l_w�s�$A�%i
-����Q��)��ݠ���;���{�p��C#;���M��Jnz�Q�T�G��ΐ�M��F����{]��Uq�:3c���w�ά�P�ܹW���{����$�0�&M�UO������l��O�ѿ���o�Py�k����'6�)n���^�5 �I���Q�r,w`�OHj�s�LP���<g���*D9���������޹��g�lcGA1K�6���v4���&+�\�+_̓|`?ҡHn�99C�z4�-д�p���4
�\B��]�Q�#��W������v8}���+���˔պ?��i7Lw�j�^s!�uwf�<�O��<����P"���ٍ��ߙ��I�'J==�'��ߘh�e���B�����m��/X"�鬜L�il!;���Um��K��t�)_���-��[ɺ�i��{NZ�'�4㇑��i�*)J�䠴�Xz��C}�3r�j����lv͒�~U�޸J�/�ZfˉN;��(g[�Ҡ�_�$�>�m�M��O �?>J$9���c΄�p蛲`�"P�F�E
��y�~(���͓d�S�818�C�Q�������!��\��� ל��-�����״G\f��nu/�$� M���h��_��AT w�� N�������)�J�>� �
�t!�T��3�����R4#���ब�D�����G\�S�*����$[��a���C�`�_��V�YX�Ŧ�zz���`��,���.�����r�ޠ�$fg>%+d={����I'���X@�M���I������@O�uV�2�¿�*�������7�M���O��{��������i���aԃ�FȈ��[u?V�n�/����%��8(�f}׌.+9i�*lY�>�*�q��u�I�����x�1�I��_��l�� y����E���W���@�f(���Y�q�Ǥp���Ĳ4��{�m��Цы�W���}��mlVD�y|�NgWB����4�&�r������3�[(8�:����oƖ:#��Pi;�]���=ո���f6���&�{4����2b��e������ċ��+�x�A���=،e�bT���S7W� AK�a?MF���썠g���(	�[���bT)8I�@5�`�_�⇿�7�͞T��������5����,O-�u���;�9#	� ?ɾ!5%s:����"���&�ӸRS���`���OɄ~�yz��j#���ez�]���߽��F[��	4������̷I&O[��B*��KS=N����Yۏn��<P�	P�%>/��ȝ�����3ϫ,g9�eiK�����6�%��|��3�;�#pvg�e(��B��a�%��8x7!��a���F<,�����Q���4(;�(�ؘ�Y
�H�7�u�m���`�d�.��p��\_�UO�r'��F� y����O5Z�%�Ȋe��r��t�b?���LA��Y�x�D����S�6^�@��d�ĕ��rv���"L�E"���o�"� μ˽K�D͂,}��,�=����W2-mǛM��d�B�j��ܛ��K�1X��#Y�dC�c��f�����;$�_�d*��C�L��7�'W�e#�y�V���cL)9��:�|KY�KB�S�V6U�ʓI4:�+. ��;%�h7^��Χ��R��A����tm�JZ/��#�Pg��B�5���~����?��\Ǿ!O���W��Z�.���f��i�
��Ibu:�U|��D��>�ސ�Ʀ�.@2B@0D[��,_"� Xs'��0P�.�����a�r���#�i�sXg�
�D���`]S|r��(����C͌��=�5�f���L[M�Ĺx�֣]�U����h`�A�w�����4-�Y��hohK�-��.�����W��
H�[xE�%zhI�H�'�tѲ�Ȯ���p�g�.��7Se�h��{!Q|,�3{kl�Cz�'�ֿ7�]q��m܃\V�I���5Rrs<:����K�y�#�.�У�.p�A�?9���͋My����[�w+�4����F�WI��Ԧȩ(+�@����e-�պ��
*R�Dm��\����J��m�K���@�_&�`o��b�:�VcX8�t[.tY�t�8�g�jr�Ɗ�i���������*0�����Z����I/�tc�#�<er�u�8�Oxe�Y�a��Q$��=�:�A��L�iϬNb��e����؞����r9+�%��Eզ0��ș�E{SJ�u�9���"HW��-�u퐵��#��L��PrE�~��=��A�`���Yo�oئ����C.#{��Y+Li,0{6�����\K��&�x�u*�K��s����?��Q�͟+(-��]�#R�T^Y�K5$P!B�$�yל�'}��3{�Gb��챽���Pջ�?�ho�<�7�^����q�q��q��3��N`a��?������v�$�A��ɒxh A9��B\Jv?���Zq�L�*z|�ץ��!�=�g�� �Rj`�v��6��Vlt��fT���ZKf���L�'���3)�V�T����y\��z�]6c�^E�Lu4��Wa�2W����y|�n�:9���[~�=��c��I>n&1/�������I���?��I���M�����]����-��9E�nD��������]"���WE�����J$�)�t1�R��j=_�N���f�D$��#-���@�S�#���J{��3���z���v�,t>��$_W�
��/�U�F�x������EkVe�7��"�e61�ͦϟ�q��ힻ�2��7�AM�K%d�,���E��l��F�:?)�sˁ�/���D����Ch+��"c���1���iб���#�Ɋ׭MdX�ׯI����Z%s]��}.��d-IJ��xY��&y^��}�qV���h�i���Q(�&�R,un(�����sܩ�$�@Z���Mӎ�SķNt�z����a�jƯOS���ѷ��u�mc�_����������m�FW�aee����`#�`8x]����{ �T�}�N�=.͞�dh�b���ap�W#e�3��`N-�62i�Ϙ9ȉFF��K�<�8D�Uo�RFljE�a�h{��qT��9�_��3'�SD�4�k&��Qt��y�%8w�����Y��P�J��f'y.W٠`����f��@��z��x`��� �y��f�̫����qR�)��� � �m�il;]�M�^�.hY�!ps�A��V$m��� 7��&�cfٯ}ޖ �-Bq�݁Z�ǭ�q�ҍ�����Z%����˛��y}�j{�ɏe�Pe�����4����:WQ���?�=��Lt�s�iD����du������ �k�&⮬W�@��x�B���g:����t�#��,�&SE�N�@{C���<�Q��+:fNB�K��u�@�z�Y��+5e�ڨ��
�_L�_�R�%���c�.��]��J}o��"�)��#��&�ic�#D���-=Dp.�1bL�`)�~Y�W/��%�%f�3&p����Ip�p>�n��40(	��V.X�!�ԟ�'����x=ƺ��<�ҟA�s�&o��?s�i\���C�Pc�S�����X��+�{���'1�f����3��w�5Z&�r�*���گD��?�s�q���c�{�nd$���t�K@��C��r�}*\c�c�K��`��xĉ�K�/m(HAC&;x_��L��d�l�\�q&c���&r?�S��ͦ�x%�5��ۮ�'#c�M�sҼ�"��I�pѨ湳�l��-�7�Y�ǺeOm�b� r{���JEJ��-��M�>3l	}�}֐�>�T�&��7B�#��"Еv�E$�������F��v��K[D�ZDMy=���8Q��^�d�a�N�\v<�G	���_�Lz�y:}C��g�O��$�,�������@Bj�s�a�V+��5���A�ܫ݂��R)�e�xl<��T��'ɻ̍J��xŭ��}�V�������P���D)�%J�.�����DZVʇ�~��}�ЪSͭ��C�����z��_r�R���&Ֆ��Qp��b����H�4�)�g���}�=t#�D��;���f=~��䩖t��w�7����eE��p8��M�P�~���mc�g�m�5���:|LH Hf
�����i~2<�0u��!G��W�_t�_��U@��UU� ���Qa�[D�o���H � �K����A�qR��d������5N9։���ɪR�t�}����R�����n�q�q�4Zu+~��I�e���	*(�te����%"W���%Z��Gc7,7z������"�A�u�o�������}�K���`�m^[�4�����U����蟬���X�Q���!��F+_ܚ1$�Z�Ц�ӵ���2�fo�}�QA@�!��JK��:p(��^M#K��S�R�(EH��Gz�����lU�$ؑ�d]��i[%t:~(�J��M�X�[�Rt�ߵYFu���Y����X�� �v�i�hq�}&t(�;`�.[Mو0n&SeK���x)�,��ќ�;�#Y!�#���қT�$B���QңzOl��Һ�LI��8��*�F�QZM�^��O������W���ө�u[үPEw�z J�*SyA͂�})H	�lU<j�u�-i5#�eCݸ�b7��K�[����\��5�fŦ��.J{����+�}%�9�j�aǌ��E��ʵ��K�qe��E��s�l��7�Fp	��!j�R�=��T�W�]��)��"ETOT��(WJ���$�����]����[ N�Ӻ5Nԏ+tn��������:�pz�mU���D@õ���F� �4i���o��J��!��Z�+H��7쒗��%D��J�aO_�	'bX#4���F��`%�u�"����슛�����7���9�[zpd����Z _� ��~�J�L0�⠴���@5��25�A'ehQ+�{֗�~�(Hl�jP���h=)*�۟jvĻ5�	�d]-���%���b��y� -t��:�N�)z�E�-0��-#R�t��Q�R
DD��QV���c�[nU)����8�G.�I��lb?Ui�G�m��~��GA/]+zL
�B,l���2wK�  ������ti�e޴��~�W���6��=l�}�kҪЂ+i�Wt� ���] ���@_h��鯺�[Zl�.ȭ��,<�j0���h��F����EU7M����!���Ҥ�,��7F�"xWܚ� ,���Cгm��J����Ep���U��G.�g�>�=�'v,\2�j�;4jL�@�m��񂸿�Z2Au�p]�tL<���Q�=�"QRJ'��tZP�D׵��+^�T�I�R;@T���-*ӟ�}���J�Q�$4$�{TU�������L�+�d/

�t��'#�
-�
���7J���R��s�eN��TrDSs�"��G�R5 d�+~9g7(�Kg�[}�s��m�j]�k�����G�S�*�L~lVq�y�ͼZ�_r��%�(HI����h��[RiD���4����Vt��mC��-6t[Q/B�iQ�>�����ڕ(tU-��֛s�N��4:�"Iת��$��Wm5�U�F� j �S��袽~���Go�M��Q� wS���uvVy q�kt�s�1V1��h^{%��KO(1&�i¾�>\�	X�����n=�4�H�c�ڱ��;F�e)�[O"�"���������v��lV�~�3JiS�N�"&���u�K����eH	T)WH��W��.�E��$ 2*�_m{B��=(��+H���vl�F�덍�����" ��uK�5���"V	��U���텘����=�E�X���򬟡g�f1"�y��r�V����r�W�=2T�wQ�e�r3� �����*�*�0�
���(t�:�EmiQIS��)-!�����DG�4���o*��}�A��G#�ׇE����|����O�HU�����i�_ڞD!�-/n��*/���5^���w�5�HG/���S��j���.���#.��a8=͛��� -�Ot1$<Qg�y��[���$�[�s�߾�j�O�I�m��-�\l����^��L�(��-�i�|�7�an��B߉�&��֌��qG7��Њn�{��t�mzq������ *�v�����Mm	u@]k�]q��K��19N�J��Q�]����zh��P�J�#���W�R5%�h�Yb/�� ��mi��&d9V�n�	i�6O��)U,��z��.;���	�e�n���r��8��$�3dd�%�����Fn%�H��4��?w��[O�=e��&���zqڮ� ;�خ�^��P��7+H�H
�J��<���6D� ���hU*�Z����/6�%��4���T�-*P҈Ui�T"ꨫ�_t�������;2��ժ�>���<Ɨ��,܃�2�>K}�gD�	&
�<'��Y2�+�1��C�5��/����-,6�\/yVH�W+Of�\�����tH�[�[���u��.]�%�/��-�84I��H�P�z������UvU���V�kc��x�����*"��.���l��)A�`����ޑKj���؅)
V�tHJ�G��D�!�j�D��%����n����s��p���>cc����-E����L�T2�ſ���Uj@���;E��ey
��	�ݺ�sT6�)���*W�<ߤ��e:�ms��S�ꢸ�E��s��?�A�		��>)]HIR��JDB��"/�U��ċ!�"#�C�DAUhv�!RG�FZR6գ0B��AE�{��]�� +]��{�F�L�E9
�܌���>�� oTMW�WU*���c����tY�A����_d��-r�z�'��7W�Q�L����B=o�t�[����7�u�m�]f�7+h��f�{�:=��Xb?�$���Q�O��HZ'MU(Et�t�&����]h���n�|��}�H������(5E�k��ϭ:� jG:�~�q�+��T�zEڪGT2eiX%��D�� K� E��l)�h�2gM��h�vEx���Q*�腄�w�P��,��n�)4��qF�:Eonڒ�ԊRb ����jE�c+g扠6�v�p�\"qN?�L��&����ǳ�zk-+�\��a���^��%R=��UF��V��� �e�'C�'�?tI�tK]�&T�'cO]7^��4.Pz��@�d$&K��Jڪ3M� /x�h@I(z-uM���E�C��V�ٷedf��X�$�6�"�"uN���XL~ʜQ�9��Adl9���z��`V��{��]�u�%�^x��p�@y�#~k��E�-\ڽ�{s8�2ˮx�Q��>��4KtЋp�\��r,��_-[P����'�D��׺��T�}��b�[���~�ޅD�Q�$(҅8��Vʑ�Z������J��ޫh��"'���#�"�~�S�vxhd��s������$�Rs�K1�8���)Z�Md��Z��d�Z�k�T'ǌK� %��O����7Rɸ�n�wHw��#��9��w����1�e.y �r��6��A������t�졪��ed7\~��)}dF�`&�Y4۶�����M�~CF�B��;���:+��v���H����$2j���E��$�/@�^�<i�-�H�;@�G�2��EJ *D��Z�um�%h� �e�4��T]�iĨ�Pn�N]���*�wn� Wh_������[��g���ɷ�䷫�Su�+l=��Lv��!b���kc\��K�-D���[Q��ds�	ݱّ�3�&/���Z�[=��ز��X��JC �M�j���f��(wN�����%qE������ ����*��U��o�'��!p+��='�RRt�)��u%�ڛ���IF���U�vD_/Z	�}`�_R�+(����Z��w�.G�=�ɭ,Yo�.��J��&� ����J�r%�ċ���|aA�=��d���~,ʲ�u<cbV��M�ۯ5o���q����r ]$��9�%Įy/>^o�ǝ'���ٮ/�A�;�L*��<�ߑ�mJ�<�)���؞�(��*uU*W~��j���TB� ��k��WbZ=ב�#ʄ��'�p�Ҫ�G��'֖@�y�d+f$��$-*����]t��籈�n8�:���uU�W��qe���}]�Vt����xl��u��qոK�pt��˙$c�K��s)�ʦ����1�3� ]�jX��2�L���ǎc�"��W?6��\Zt�ump�inc�*�!J߆�	 ��Q�}�T�;N9��$puNѫ`ݲ�.�@���C]�b�}�v����=�ْ�Ӌ�$�֕�4�ZT�צ�;��ס��ywBj��ԫ�����=�*�Q	%9���Y�~7\�⹇��Z�7ӏ��۰�'9?6O�ڼ��̰� �}�ge��Q#\$\\�F%�6!b�"Ҵ<�3�)�+t�o�HJ�� �=k��(��|�{li��� n^@*x�qUj�ǹ]nҮ��h��뤀o�6���)��k��I��z*з�����.�W�T5�H��(�/bP���}������+�V�
2E�
�wU���wWb�G�z���@�I����:濅��u�f\gbyS�Z�`���[a�v��������ZU�5Z���1��-8��ʤrQ	ťstۚ^���Q���=����{��捴ZO�T��"���PSI�R�t���R�yi۰������TT_u��(d��MAE�W���Ж��<t�����q�%�<�+K�A��9x�O4s�
8�y#:� ����׺a�qƔ[<<��Qo����~��FrM~L�4������w��|���lO��5��}�Cd㮗`p���N�F��]/q�:�s؇�TARJ$�5#�PE�� �� ��%)�~ʝ��ou�k{���P���"y�UŭuF� D�ǜ*k&A ����>������qǮJ�w����-'��mz���]�����c����K�7eß��F�wE��3?�z��$;" }C�|c(�
��/�GCHE:Я�t-�.+��a�O���*��.�үe��O����6ޗ�`ۊ�B��;'R���ivF����tsg�/��h�)�0�#T��a�cM���ޓr��jk��-�em� G9#���� 4�1��g�U��%�C�Du� :�6hn\5���\:;#�B��2U���8gou^m�o����n�8n�����7c�� ���Hu��S�����U;mM��v�{�tD�4c�\A"�Q.�v��N4"_Je_JM׈u�.����R�U�B���xU��]*0 J=hL���v�:����U��^>�AIڶH���g]d���b�ĕ�!�c��f�'|<�x��C~ȸ�,��Mz���Q��S�	q��7c.����}��m��/�<�ڍÏ���?qzV/��pX����Y�o�_ʼ�h��'!A��_��f`�8��[v�7D��J��k���M�گ#tjK_P�=�S~ؤ����j�^N��!N2�/I9���!c� Ů����W�(J2��J��D��ӚDB�����r$��l�4��Q5@E!of�AW=nߋo�	����'$��,�K�D���a�\�t���^1����(c)���\�w���"����$X�s��<��(ܲ �>�Ξ��G�F#6�"�
u�� �˭�Qf.1q��s���ڿ�x�!��6V<8͘\�����di�5F�B��BT�a^�I)7�RZt�[�*
�k{����z�rQeΕ!�J'4��Ү��Q6���괞tTY�	�1|����R�)A(���_&��UVϲ�u�/Zi튻R��6�m�͎�˽id��i
���1�_N�d�[yj�e���_�GЄ���X_aʳ'S'��h��ǋ�,�Үp�q�^ݍ���-��o�n�.x���y�����z���|��l���e�\K�S1�#hr��f	E6	�v��U��t��]���+��Uh֕	h�P�F�WQ�&��E"Du�_e�^v��)V�*�Rsu����u!�{l�Hd�pWa[-��3R�M�:���A����ʈrN��*a�S/�XUը���!�[��;�lp�������}$L��-~k��Q�;�d���0\M�^l�%
��ū�a����9��.}?�Cr�.O�Svx,��\����� ��9�<o~����/E�DJ���_�5Z�HR�K��ڡ�]DP��3o�m�{�n����d7GH_i}�	��}��^Dn7j��COz��{�J5T9�H�_��{^�+�t��?dRDa���c����<�ۅ�A�X/���nK�\%rM�D8�.n���	�P(y�bs�8q�`�Ņ��Z��c�i��<�#�R>�}Ku�d���J�J�<�/X�x]��i�O)�W�(���*㷔s��A�1��X��hq��4���jE�S�-��g���Q��V�+��.9-�V;l��d�`q����?�e��et��*�!�p�#8����Ol_�^Ɔ�{Զ͓	-Q/v̩�CTޒ�u@DPJҭ!��~�~�PM�h=�g�6��r0WB��D@�� x�?��%Rn��Wf��0ќ���6��'dW�� (��&��+�!�.
��4o��i*�H�E�����_�7��I�!����GC�C��p�.q��[�����4�3�����/�n;*�T�������.9_��~�����Ǜ/��nU��qʧ�����S�P��G�+�P㤥���D�ʯ��ǵ��q�� ��5��;�+�L�t����IA�k n��ㇴ#�� $|{�$3��W�-n�x&C��âJ�}ߺ)�|�DJ����v���U���El�ծ��#����M��r��2�L%���كI�U'�sZk�\Q�YmJ����Ӆ�F�� �{�lYYg��~x_8)�C�0��r�U�B������/�4H��^`���י���G��=n�ے15Rſ����j���+�dki�2GY�*p݁��� �� ��c�Mq.2�7�_2�q6�gĸ�o���D�li���XՋ���� ��� D  !1AQaq"2����B���R�br#���3�� 0CS���Pcs�� ?nZ��T��t��pE��m!9��[YNk��N�	�vYk�����S%5�w��ӄ�Q�����T�S�Jj�U.�T٩���voT�C����H����,�����x��e⺺P�Q�4���uW��arT�U|#�|>���[�� �,��S9$O�\VC=� Nc (��aDǪh�y��f�% �RdV��a2F��a!>^)ͦ��`�~��D��S+�@9@^S�V�9���u�1��Z�tr���h�_XԄkg�����9��3;!��:�Dh�I�cI�Ȣ��#�DUT
h���7��@��m�PaӘ����MokO찚�Đ[�)��e$땂=Q���K��6}e��2;�ki��Y��Hl:K{^u�:&����>�At�yh���L���z��3Fbo1�.hh.�lx~]��0��?���8��� x{��V�Z��&m��f(E8}��e�m�m�s�A�0�ߺ�>c/��=�/��� �=S塅����1�5�):���P#��	u����F����nl>9�����1;�LH�}V�Ff�ͽ���;1i6lҋ�ӝ��)?U�W� h����� �� ���c��o�ba�!-�d��T��#�9��O�1� -�F����0��N�خ����D᲎m�M�E�`@"�;d� �,�tfS� �
��i��������M���ng�M|
.���Ϛ�� ���� *������x� �X�K�%Әr44��|Z:���FX��E�>V�48Mܼ�$'��%���˺�I��o%p�e��V���y+V��B+�p|M(Q� ���+�M�_��tT�p^ZNo��f���R�r�2�Ҁ���V~�a�ZL��^U���=���,���߆F�h5�,���Ua�N b7�A�8���di���AnR3x�a�fx���Y$�� Oe�"9��e������iE�����V �q�8}���#�lv� �j����=���E�7O �;@�S%�~� ߲&M>TDڼ��:�d�ağĎH�������&��x#9�"�t �0W��6C.o�Xk�S��?U�:}��'S4j�>i�p����(Nfrf�][c�y"6h>E������?D�Iw+�=�"��38��"s
�SNSAE�m�r��w����1���ӊ�D�9���_�&_��
���Z�2�;�ub�mD�y4�N��J-#j쀐�qT�iI�}���tf6�w�`,L����Y?��h�F�� �Q	Xe��� �})�}�\�.��U�S��� ����SZ:�Mŗh��ڧ4�.(u�P��\<F���x��5� �絝�S�'9�ӳ���Ǌ�rp�N��%aK���ߍ���\'1��.!�7Q����������Β>���?�se��ߚ���k�FT&a�EK��;�N�U%��'�OY��ЮE�-Y$�4E���L��*L��<̟�`�×���MS�RF��ʞK7�����h �G(v�&�T)<��M�a�:x&��*d'�'�f�{�]� f�߷� %�[�|kEP �����4�[��r)&��4
(-e�7o4�7��oY��'�E���~��,���~�͜6����a�N'6W� b<SI�C�C�V'������N5���ӱ[Ԭ�%u��Q�5�y���7�$q��5�<�A��sJ�qOy�n#�j���Tܚ�?�h;����vNXf�ea�5o�ܠΖQ�I.�X,���O��@M��x�ڰ�~��ěPךlb;ӲM�A�`h��I�\��ā�G�?v�,Ӑ��g���D��:�ˇ��p$�	���&]����c��u� d����Y��حn��x}��t�9��	�A�D�e�,n�C[�l&ѦQ��"6E�vߊ�빦�1�,�7��t�"����%�ou@�u��J�L\�q�L��싕mƓ�E��bS�5��a<�����e.h��8o��Z6�_È8�c�G
�D�U�]�c�
����}u	��1�k�>� �A��?�%|Ʉ]�.+��}����f[�І&`�2�o�EӞ�w���tN� �;&88L��(b=��H�ew�?�:H-��{��r�Y�v���`��mf�gsˉߕOi҄/�l���M`ohKG���Q�2ֺ�����X�&+$��	&{'Ot�#4��4	��$m0b���`ñ0�)�`� +������k�sGد�3�w>KuC� x��Q:���'�6nj��gx-�<Td��m�Y�)�"drB�d�dW�O!���դn���2��w�D��-؍�����ƅu��L[�f��w�|VY���hLp�W�s�b0,w�����>U��XPO#�[A_���4�����{r�+��?T�y�CH�i����k�`u{:�E=Qn,��m=WUC	&�[�][�C|��)�t��b�\���"8�=�&�b�')�[�%,P���_�e �k���\g,G0�$�;'��OvFe��d;Ls�?t{&�O�M���� {��#ĕ��b�P!�:L��7�E��:y�怱�#D�܍=�k{�#.�O=���͌g�owP��Px{�AӘ��[�=Vgi��˴9����a���~%��;6�/℻�����2��Qۣ�(77��U&6�>���Ui�KK��X�@o�Ou;3{�
��}Uk>H {�M�#�=R挳z�G���'�v�Hv�	��m�T���nI�7!�l�'�T١��a�\�t[��wz ��V�3���5�iw�`��#L���q�A ���.�08!�k�Xi�u�X�K����{SBwX��#������isb���i��.p����j��k�=��q��6@��.��X���kr��3N��;N���亮̖��2��<49� ��y�E��P�cX�Lq.sH�Si������vrI��[TDY���Y��f�!��g7� �i'�@�&�ule��8LwxJ�;��E�;[ N��a��]�yQ�X7��$��ڢ�A���>h�|S��<j��#����/<.&w�z��2�io��OuI�4��q:M�uM:&��$�Q��4�Rq"~�P����i���^Gu���ٲvnɏ4����D��p���B3��z2��i���ah��Gt���F����rN�rL3���o�27�� �6 ����:�����������9���>@ �m�����G�x:Ea<vI�{��`� ��[��U3��h�ӂw�e&����ȃ��H�#�۠��b�ж%uy]jUb���� �E�O��&�Z)�XC(s��|�}~ɹ[��˃�Y�6<V_����.�Z o�@S�~���3�|���@]K_'8li7][g�\��D��h�S�Z,3u��\2��
�)4�XN�!�.@�Ih�f��ߝ�<I_��r����A0�A���	�{J.�eo5�vVx��T���x�:��Mxlk�N��De��L���'��s~�� Px����JT_�i���b0��� o�e�����~�Ԟ@����S��� �N���)��X]�� H�DOvi�i-9���H-�Dv�\tY��k�`܏/r�D;(�"#��$4��ߘ�{��o\��1NK	�pF8~%�����x��0���b5�y,g�,QV�L�S��L��Nqܢ����tv\�wR\�x�H�L\�sK]�WE�,�~��	�n%jH���a�*����3T,�̢e�����0�� �4��a;}j�R�=� ��c�r)Ƃ�O��O%�u�>����>���Mj�P0�Ve9���樁� �g艀����@'(mkDp���7dq'��7�SO4�V�����Lgi:ID���^��9��3�J�2�s-�(%�h%bW��ֵ�]awi� &�1;G'�\��ˬ��� �'b8��'�`�6� q�}�i!��@�������~kj!�� <N�~�_E�~�I���0�,\G 5�eq����u5X�i M}wI� N�}ea�0������L��<�]�;꿊� �)�O�8Y��~��W�/☯��h9H��cVK��L�m�w�Kk'r����U��� $�M��( ��05ך{L��A��Lx�be�m��N���͝���c2`b�M��i3��u��8����X��t�6b��+{{#�~��x��O����k��$�q0�s�M�c���p�7�>D���a�� PtGL�5�[y�:Ja��j�e� �=v����<�3&	o�ޫ<� �����3-����bbK��l��!����.P�LЬ���hA�ߪz /����V Ll7I;��H��v��ĴvZ.�(i��%�+�,ڻ ֶI��: �k�We؂O���;U�ɅƺS�k{,�,�t  �����S1T��&2I1cr�Y!�����X�z�;���d}e��D�v6�wR,N��6�
Z���}���	�x�9�����L}Sr �4��<�-�;�e 8�܋.�*J������Z �G�7��?H��v�B{T�x\��Ni���M�.d�@#�YE�)ʩ�>F��,�.����t����o{&��&��D������EcNcnd�{EAil';1�F�Kc��<=�$:��Mq�ǻ�=̣�Jp0��((9��@T˼|�ܧ{���Dl���ñ+ �a}���c*mT&�~� o~�I2�r�V#Cd�LY@�\N� �#�Ƞ�0n�7qk�S:69'H��!O�����h�v�����~�k�4ڟ~����-{Ɵ��Ėװ�O�9�fW?I�VW��8����� w�}�W_|�#��925����u�i6�/��m#�Xj��ژ�����n�ygZW�j����i?��|��S{�l8,��sC�Ϊhh�P�Ѡ	�eR�=\�� ��0�����^@ː�Ӈ8�#��	,���<�G���♍=���Y�6�A��$R�]��"y���c�]��#�P��ӣ�Կ(�蝊0�\�z��_�2���WX��&��m�Pԡ�X�w�8������p�-:M��cg;B�����a� HY�p����w\��@�����|��5��7�w����o�?��O���E����YF����J�dR�a��F\R�D{o4��80ܭ�� �I�DC��w������3�CEܱ7� 2�zI3:���A�G̢L�R�,t]eGDh(�2�v��ߪ"%a��mf	�,C/>^_��i/t"9Wa�X���jn�����Gߗ���ŌS��8Ko�Haȗu y��C�N&�|�� ����^wOl5�:ǚi|<���/{�i�K���:}�&I�_�+�h�CiN$��+�u�j�=SG��� �$�X�+���i�u���n�K5��4>��c�\Mu��f��R��;�}�#�~����������ǖOg�#N|RKb�����1o( �>�d���DY*D��x�3�˗�@uS��=VL����e��D��ǂ��v��U"����4w�hi�Nh�ô���S�Y�P�M#� tx�"�P��(�M�ꉋ|�?o��1`���:��P�"�Q�f.3i�p����z�"{%Ϋ���Y���5��IӚ��\�t
Ɉ�U�b&�1�ܮm"�iu�2K@}?���,�1!��_�Ϙea��q)��RK�Mr�O�����p�44����(��5��+I',�u��ks2i&o����9���1%��:��G��y��/dMyHL8O�ܺa��.?�|��k�ip���� +�̺�5�mC�,[-!�R�.���7&����>�f��|F-Ak`Z�~����lns}������(t�'��V��<z)�P�,�+'��` �z�	�j��#5QĘK��
��R32��������mn��=�y#�%�@���k���  �z�oy8LAL�@&S�*G��cⵂ<'�C���ɭnV�8����.}�0���Ι��t����CE2����9K���p���@7���k�X;-���uN�j��Mk��.ֳ�V9�A���d�L���0��T��|Cv> ���t��}�ss�Z̉o?���4Rq)+ef��e�m�߮�Y��Kv�}T>)�7q���NÝX9}0��qsi0��y!INR����:	����,�q�e����x�>�[a6i��)���a�8i.i1k�T'9�#a���iAQ���&�����G�`"d���= ���x����]z"SGAs���av$����|�5�F��EW��>�U�wX��( �u���ly�]L��Mg���i��Z�B
s�D�o=�9C�*F�q���3��4E�48_S�-���(<S~!���3泹䘒���
��8�`����-qn$Ǧ��V;1�;l3�[��V/�
M�������\��n��o@�P�����DV�H�G���N�F��~|��F�]t71'`H�Z���~=�v������q10���������Y2�ș&iTL (��,LN���ԙ11�j�� �~gq����wk��n��Zi&ו�q0˛՞C�gu������(G�����N�3X��ɍ���͕�^��nB0�Lt*DO�E�;,���<���@�'��PO%^*�ͮ�~°_e�Q�tA��M:+��@$��|wU��g� �o�LC���wG�o���a�mI��5�{�KO��l�˗�N2��u���i٦�(���<�#^{m�X؍����k�9Z��1m�X� ĘO��"���ZRm#�����t-��-��0���A�����{��)kEf���ߞ'�|CLS����a�`�g��i�f~l�1�!5Ǳ�� "��1��2��4����U�e�dL�J��oĊ�+�ӡ�X�n��ټyQ?��NGa49��a�F��h$�0�q��a9�� ���#�|W�7��p����#�z/�������L��r��X�u(���8/sZ��ۗ�6�⸦�C���?`�>-����i�cI �}��g] �3j�<�/ĳ3"c�\�u4��7��_N��Gzw�1����ӗ���Q_	ԅ�� �(� aJ�tL��(�F�tL(�H(T�)R�4m�+Sˡ���� }��+0�f�鮩�G5$X������Su��$�<�� ���X��Mh>����i_����5�E�5���U�-����_c�N��g���]�Gj��h��D/��0/�G���+��b����<��	Ï�ߥ������)4�p��|\��/�wa�v�����O�a��͙��	�㶫��]�5ZCH�}����c8/��)���u�S����@��l`h�+ò��� Ġִ���6��1��H���.�U_[�7{1h�)��Lj
���)v�f<Vs�pMq@�E�:��$�,��R���-$�hSH>6Cc��!Z�,�T�CMa��R�	���'՘�$ @$ B���ST��$lc�b�9ƫ�a���wاA�x�_�����_	��[w�X��CZ'�.��G�	{���c2�+����_9X8�1�_�E�9�_/�k�������g����9��*�lO%��� ]N�y,0�7D�z�x�D�d�_?� �c���lWvc.��vU_ �k��~��E�X}�}��T�SZy��gnA�S�Xx`R����N����)�-nT��>6G�ی+_��4��A��V���we<�߰�&A����� ���� +g连ĦX� ���~?w�w6��?�1��ɡ;���-Ý�����؄KF�~?~+�����}�E���8����k�&��:Z��=�-t�+�2�^`�1z� ��D�]H328��Y�8��L���w�?��ho�3����Sc�<�G�=�-��(�ڐi���g�ɖEo	��0�D�8M�����C����&�,0֎���a� ;Z|$�LW����4�k���]k���h�����s�ֵ�����ˌ�05��?� w���$�W>�CN�����D6�I�J����n$��a�{ G�r��v)Ɛ`���cM��������̝V.w�6�5����@Q{���`�1\�Y���X�!�h�k� ���a�0̒m�cRK8���O�k��ϗO�Md�e���� ���{�u���9�sD�G�{���;xn3�Y�晁�״� � ?� H|36$nY���\(q�'�|�L�NcC�)���]�_=�2� X>��ȇ;$��9��_��@��;r1��M�l,1۞��'�t� �����V�NW��_�b�3���'�%́���ŷ�'�!��(<o�=�]?�A��3�TBrs����x����-<W$_���
s��RM�d��C��Z[��沂)tƗ]?	�-�+��5���4�`J"��T�c�ߚ��^M�F��*.��k�h�;/bDL�S��)��h�wN�r���e���h��g�1T\��ǎ��X���Yfk�b����T�ॢ�B.�q�uX��\&@j[.���lZ��X����P#�V���V�����FÚ&-����.`�6�8m��v�S�$4wǚ!��v���#1�M�'Ѐ�>c�h�F$�?��+���7�=cA��1�fg6�W��3	�s��N�Q�M�a�\�t ������L	t��sA�"<꺷@�^�B���S�T� ���(�7.���Px��+��d4�MVQ�54캓���1�LwP`����6Pj-���ǚk@����wBw�7R���+�.�\#�)� 5�`��[^�F$���6�p��z����3����0���P���g 迪.�Jn	:.�uj��4G�r�M�{k'�vh�#�5�_ˁj#��f��XC{��.蓗�T0	ຂ\Ѳ8���Dh��ħa4��x�W�.��|��X $�g4���c�HP{��M��DH�Q-j�=Jk{+1J��.J�֬Q%f�v�PE[�R�����?z�s�������}]O^ϭ�缚囯��������B"e��ihàf���q�����=@SF��m��ĝT��!r�:E�"��,n����=~��"'�\�s��p��I���bԮ5�vz0/�C�U���A�pv��}��jv�{ą��׍y�~�X<���H���[�;EN��x��<���s�:�\.�U�*N	t�A(�yu�y��⟟w�2��1�De�QX�S�_�p�-}�!�&�;�#��E�t���
�j�����$.�ê]DV�@�s�Rns|��K�d0�"�`f6!��ןS���t!���z��X��}R�궻]V�}W#]d�W!ԗ�d�M�FN����?3��YA�\"�J�K�Ӣ|4��Qv����3�fa{��:t��5N��;l�� \	�T.��4u��Q��0e�N�d��-lF{[&�#c�GT�� �ҕB�fJ�I�S��'�>]Z�OG�E�����m�Dt��G��bz�5\Sy;K�ƿ0Y{Z��z���M����\��='.�1G�P=�������q�HXS�V�*Tq-� K��"p(ۖ�*��@�љ35����C���L0�i�;�,ގc���ob��P�E�GD=����`�}LG���d8Ռ�������I��������F�3�Ylb�Pچ�4�7�o��XSu�%T�����ڋЦφ�3�J'z�O$;��ݏ�[���^܂�0O�؏^S�a�_�ŧ�`�J��#�2��v��E�}R��c΃֊<���="�j�YR��tp��� {$N�[������U�0�g��@n�%��[������>�&��W�p@�.� ��'�|���iW��d�;\5�&�����['~׎�<]t���O�����߇	߷T����\�> gU+Y�+�E*u
'\adڿ�U4ӹ�D��Y�.1����_�R�D�OH���O�e�E�>k�[i�	�{���Ww��:o\4en�-coS��<@�����vgK�q�v��l=NM��݉�u߰���ݐG)��с��R���^"���%l)��qӯĠ{>����?7�@��0l6��K�\8ap���
�B*�:b�����l*��z��]�K�LG	9ۘ�j	\}�t�i�����O�OV�f"��`���/�.NN�H�h?���R!��ulePC���|VW�
jcS�93��h*�7r��	P����i�}�Nu���;Ǔ��hc�T���^T�-�k �EV���Č�̈́�8�@�� �H!S܎0^W���A4�ʩ u�P_. Q:�b{��"7�����z�W8��O�k���Q�cKSݵ����o��?̂�h��=$NS� ��o˼��J+-�Jy�."Ĥ�T��T)Q���p�]�j�P*�T
�Y!6�G�6_��s�=`�n(��IO��L��s��1ZD�X�G;m|��:���nxZ�1�D�-`�dَK%+�%���J	~'C�m
$�kC��H��Wެ���
o��B<��������9�y���d�Ѯx߼���	�.=ГT˶>�_�#�y��������"p�T��htEL��vQ/RJw�L�f)��l�*�Z##����_O�n~gk�~�/i�o�hCE\�b�0����ye~�F^TÅ�ʫB�f�u����r���b��w���4Z�.n�ɰ����R�P�j�-xx�#��G��	x������,�6��GTK���ˀ��Z���%�EWcI�P�/p���)D�q	ø�z����]G�&��J�n�u=V�\�>)3����VN�W�;E2c�m�횾j~,!H�U�veԲ-�� ��Vp���z�����8B0Jf�������,�s}�J���R���,�;o��.�4��������Nf�!ˁ�@-�	�w, �΀�C��:uܲ�c͜�\��A�ޝp��r����:#+�`�e�����b�t\��d��</j`�Q?-kXmxF�p��x��j+m'���A��WV(8�����lñ�~O7J�>���?��|Ԣ&\�F��5`��j8��$֦��!׉�нԗilᨧz�:풝��
���Z�K�?C7K���K����]Q�d��^b��(�/��L���>_��`��l�tf	`�zө�lP�4���5��7}?3P�ةJ�T3���ξ���5��^�������Z͎�� ֩Ρ�䩡�\�Na#aj"�'���ei��?�l	rb��L�ZM�����쇥�fe�,9	u�,R�e�ڔUw�&N\Q5�"����S��{�� ���ٌL(�K6˅nm#���Hܧi-���ܝ�ʝ��!��#��Lʄ��丛�Ӣ4�`[n=��ݰ�^��F�������.��^l����9]*����qf�����#� b��y"�N�zjg�7�?�S��W���{�{3���%խ��9^0�)��h�LJ���w�`�C����P�G�E"�
�t��'��G��	"�;�'��f������(
 �<[0d�T��ׯ9[�Ί�7��>�`�C����b5٪%tZ�BQ��^�8W��T%rEʬd�_�9�˕
��g�. �3^�W��l�|6+G�9��LJ5B�~�z����T&�7g90��Hh{h^Y�tE�	I�bW�{2��!�[@�{¶A��OiN���{2���ԑ<�X��$*��%�\�JE���ú�'"u�C��Oհ2"Ð4]*��OR��B���f݀�tIy�:�32���v(˟�Ƨy�XG�7BtEuj��	L��̀�D�Ϥ.#~�Z�������1�-��6�ǒ��+��5+ūS2��_�η�.R2s4 V0舌�IT2��mk�%%�t�(Ed����\b@���[�S�E8�[��B��(S��[E]��@R^�Bn��/u,֎��tii��+�����D)��l�_�c��.랫?0W�wx�\��:�mך˽��^3j��ɑ~ ��W�C�ϛG��0��ߠ�Z8tR�~"x�͍��yk)a�8�f7�1�+'�ʣ:��?�Q������+� �N{�:�^ϔ3?�̔Ɨ;m�l_��Eg�ł3�o*�P6�ʯ�����V�(#��N��b�R�	<"��Q/�Tt[Q�
���J�ӝ!���'�{Y6�h\�=$����db�&^�؉��"ѐ��<���XW�R�MP���&�z���J=�bA������ŷ�,�'zk�p�-�� ވ��n�C�؅`g5&�jsjǷ4��hǌj�}��'�ώ>���'���x� ������~���8�4�S�s��v�1'�Z��B�S� �F�������!^4�5g�("DЪ��WX)D�����t6�K��D$����M�܄ܰMEbgե��J�MjZ����Z���">P�+Bh�D��6����_�c��nJ���P��Ҕp႘���~��;��W@瘚��i��4g�X;RѾ��"������4��F�K㴭Q7���ƅ%T�Y&v!��dAa�_���ւ���ĠQ�[zŦM:���?�'��敖s>g�)��0�Ug�`�0�8Z��b�0+2�ŒX�w\XV*{�t��7	�-���X�b��?�� J��.ʎ���9s�Z�����kQ4k={	H�I[c�ů���?h��N鮎G�n�;���Ќ�1v�K�S��.Bd�b%����^7Vu��D"|5m9�ٴ.p��F�W��8���/5�!��0_�D#d�(��ϩ�}����&>F�S�-�,DnB�<���w�V�[�#>Y�|�c{	�פ����2��Q��JilZ���M��T�P��93 ������,�Lj1.�S�UTH)����������m?�q����۪1O!�i/���А�m�O�Doa�&	޳y]������&x��x2�.�"W����Q�Y�QI�V�-��ɾ�ri�"3�Z Xg�.(5r=��B���2;-�Kc�2�"z�ԍ��I���9��
�cM�FW4�j]Ѣ�����wd��k~נf�|:$��E!i��M2�J�bF�f�"�yT�^��:?�����<, ��RXa��b��En�.Z@ �P�b�eB8 H]V| 8�Q�_��������s�FU�9�{�����?|[�i�S#d%׊���g�x��^�%&�"���Q�{�����-VAE�<�W.Wq-��Z+!�����_��w��q��G=��_�c%��0Ir}K5�޳F����tiw7���7ſu��<�(8zf/A4�ԡ�B����.����Da�%�xS�D8��7�8�N��E����
����*e��lMJԅ}�����	�r�7�kNL�G1��
��p��֟W�Dv�p����W ���}� �Hp�0�FoƱ�dL[�T�U�ĩ��+KE��k��I�;��)�v�TT�� n�����E������5 /��Oob��!^d�V���K�n�֡������]��%�� ���Np�g���uuZ�7�WZ��l_Ylq�b��=³��U�j�$�J�����쮬9%��|��J�1��?[�M￥�Թ���+��x����Y3f��!���ي���G��Y[�Ҁ:���r�+@Dc�m�R���`�sm�_��V����LNN���e�M�poa��W�!P�8�3JU0��G/zT�6#�E����7�� ��p&(J/�EX����4B��PS��D�H
��D�u�s���3���f`�ve�Lϩҋ9ӆ��ځ-:@��-Ւ!'�"H�:��ل�D>Q2��I<B�0x�n�(=�2)���
�%�Y�D��-�x��������6����>e��6`�;	���y�M����h	�Ȃe��I��Sҁp��Cx��Q�r��"�d�A���_�Ҥ!�ov��եO~#'���	¤~���� �oń��xzP�Vw�HX���ShҕHc��*���\�r�~ҏUq����>�!ҕ��@��mޮ'��n|jei,k��)=I	�S�˙�c6�ؐ�e���ά����7@+z���1��mZ��!Ф%I����)�GjrBP8���� ��2R���\�,�&%mM�i�� 
|�A�-��/��|bS�D���V�崳��}yP����DιM�!zXf>�[�1�����Ƃ���*�㋧>�J*��2>A�q7�
��Xy��y;��n�H��sK���r���|�TF�WYB
K;�ڥ�nֽ�ֲX�r��Í�fp�x����+�ZD�z���H�4,�ǴI�5Q7��M#ƅI-�ۧV�;�]��.Sm>��xs�Gn��,��Ͷ�����D:�_ �������EKV���y$�Dj�nU�C�#��P+����-��ׅ�"A�gfJ7���DZ�r�"+�4<��GYo��7��P������J]����2�ff��; �&}A���QR��a�8�;��"���m�<�7�C=�d0UB��J��vN�h�_<�@k/]����xf��zeMy��ZA.���N�-Si*��[u�L�~!|m6�@0�'x'a�UhH��J��(���ZN_	5�@�n��olI��|<$ȋ�XJ���]�&����ޕ�д�I���R��o`���=>C
�����П1hO~u�az AM7%��4��+hzK}�nc�@7im+�S��m��lc�B�cH�C�w���,�����ڲ��&�^��#	�I�ʂ��@ 1�H��P?0G���qI,���B=1�)�a9V��O���8�(���N)A�W�vG���o�bd6�
Y���z��Z,ML���ߝ���̢��V�Φv��}8u���<Tp�!"ci� ��oI}V��n�p��'�lPݹ��_0�J{��lIZ7S��9��3x�2���K��T���-�*��I����d4��yB����N�0�JO�G�3+�Br�R���@������g��%�g{����j�W�8�P�sZ[��\�)�p�T���pJ%��P�3�^�6y��8M(L;��D�Y��qZ�pW~(��]>6;�Uty�ӵ�)ʤ邽�f�(�	�>��� ��YH�)�}��IB����e7fsF�g]aL9+[l�'j�j�j��IRo�g����U��-2�7���@Vrȯ��|�G5"œl��Gg�#͉\��Gm���fu���rl5��X�.˛�΅�4L��|ӫ{�H���'ѩ��\�	#3M&����*/@2�.��m�"��Y���8�����f�Ϟ<R|C2<8�"wcC��x�FN��$3��������*Kd���ENV�E�e-��Td��ƞk4B��F[j̢k�Ԍ~L����#Gv�)֣�I7*������z˓`�*�Q���,������������:����7�Ճ��q+���ޖ+d�m)�O���L3T�|�OիƵ�����L�mX�+������`u<���< ͣSu�D��Wf�M���4�����~�('N"�s���U���Z�/�*Ҕ.J��зoSۉWH9����(3��:D�i⤓�@DHf�W*`�P��S�<7�o����T^D����nvV3�rğ�@�A��<U�t�j^��H�U��n�<VwC��V�?�xm�@�,#r�&�2@3I��%Hd�莡t��7�ڄc��RPw3u�ׂ+	�Q�/%Fk(��Lԝ��$I]��YRU���M���Tp�P�/X���.��3�?��r���3f�'�'e�I>%�׀��w��&��"�AG؄�
��+��Gr���6k�� :�BYk���fO\�3�j���)�/�dГ�ڋH�T6�)���j&�3�KTNqyQ��A(�m��'��(����h�
d�� A�8+a��[B�:�S�딈���E߮�w"S88B��|R��j1W�v��hi|����C�B�7��.��,�Q�5����2�R�R�젂�X��Hy�.B�%�fܔ���A��!\�MH�E��AZ�~;�*q68�+d %` ����Qi�7K�#�r|"ZZD�����$�_�P�5������8������v�4���|紁��B]�
������O����4��	�Ys5��~!�>��,<,�̂" y��㷓�{[8��B�R���U��FX|�)�JiQi��y�]��Ȋ��b�z�<Au����),�oJ��E�J)Tn{����@X�
$������˼�bk�p���e?Ӣ'-عg��c	ń8(*9�H��>�c�do��F�h�Lri�悠��_M�HQО�����K�9��VobrGt��^�:����@s��dO?����8�x�+�v��D�L:�'�`�8ѱ�&\{��4Ը���-�mhP-� {��z�U�U��#�@0�S�6��O���]Y��{(&<UH���`��;�#x4�<�!;�d�q���Ez�
�"�=��a�e�0�|�����A��@m��=?�O4R�[�3ߖnz��fL�4z�&�N�����!xu�҃-1���ԣ�9��{U�ѽE�r�er���"E��,j+i�%cЧ<��-�[n��H��39���1����ޱE�fk%�y�w�Dtd4��Ƿ�Y<���o%�Y�m�T��m�b�=r�]D�{�T��7�����s�u���EϷy��pC�g���.��Tn�543�J2fa���Yy�c�5���������,|@L*�n� ��7���7!�0nQĒ�!���@��*�;R`A~�K��Q7X��e��f)ځ����D*J0����)�U�1�{�lk�(��!6Mj�&�Ѓz�E}���=�HxG{�N�zcѲ�|�\6G�LG���F��b��q�N�5�)��=��$b/Ļp�{�{x�k����w���������x��}Ky���? �$��?����W�&��×<�t�� ק:�|='4���ޠ�o�v���_�*L�JxR8AZ�	�)��8fs[9�Ԩ 1QY�hqPƜ�u�H�ҡCVɶCx-���V�B4������B�O�q�5��7BrG�8uZ1SAq�!���D[U�\�1p�K��B�����]�]�-9t۹��T�_HJX_�4�\��~z�p���JX�@h�d����0��l�zQ�,��_���$���!M����M=��y�^`7o��ʀds�v�}U�d'�B`񠌤�*z�'���տ�.󨶅C4�b�{�@&�h���M<�+~
�2�4��>7�E��Y8�O
�eK���e��B�R��.�+���;-_;���_6���1�h������:� ҈ �c?�GR�wx(�
>.��V���o���>^F+�%�b��֐���l˕=����~���l�>�PJ����[7�ha��7�߀]cS��ڱ	h�y��R%�:zI�� �h�t�����S}�ځV$d��5��Ł�zغ��d��0���ې�Fۿx6�aZ��p�!��^0q�F�c$��/J=���*%��$4K���Ro���������6�Gz��&��k;���ӣWty��粝�"�,�
��d�_-�u	��}��jd���]���@.M�g��]���n<���1��=Y}l�u��+���.�.�/r��>]�n^�}���߻?�w*��E�������˖��]����Fm����o�};.�{x�L3�fkػ��_���^�D��JO�>��^�Q�,~bpe}'er����l�F����/jF��!��n��?�|���٭�g��7^��X���v'f����?]c[�3ߓ����b �=v�1��>M_�j��6H�~y�~�fi���R-�^�ِ�JfsR%�V�)�:���'=��z��\��t&�֓��Q��F����x�aҺG��u,��Z�iy�)�2E`i��Ø�o�}��1\&C_�� ���z�S�}r ӫF�РJI9	��m��1�K&u@x	@�%��m�3�y�C�����?@'=;u 2�T=�,�;�@��ԝб�u9,8Tsp<�gp�a!�,-z]R�_���)a϶J�P�Y��؍�70�? 5-555�@*!6yj����!yh���U�'�"���9A�-ET�7�;�����P82x���Qy(�G�9����;�E�1j-'�_e�����m����CK�,����z&��Lݷ�z�-��,��}��lI��?N��nd>Tт|��LAN^�3N���Շ���	��o�[ʋ��ùM��jM��Q¸� I�=��M��)b����?� �zw�Y,�*K�r��+k�L�jk�P����	�Yg7�Do��fߠxL��g�m ���V����+ҁ�����T(�t_��������D�:{�L�5$��^���Ƹa"}D����3��"5���=!"]��C�z�3��ՍG�k����]������e0��B�xf@�&V���sv���Gp��:����W�e~r-k��w/(Q�}���5T����|ЛrP�0ȿ�F�3��+�ЫlS	��W�0��PF�k䯱�4(������UӥI����Nl �ѯ�!��xY�g���:X��E|�����c�Ԭ��$M�!oD׹Ð9\?�_8�l��f��/�E%���|e�U4|1�ߢ�N0�P�1X�F�f�\�j���5di1z��ao����߼��R���A�'�_�u����)S̖�oױv4��w�ly�0����Q8X/�4'U�F�]o�eS����M�W�!�@���I�� ]��~�1�xdk^;��h~��8�]����(?�Ƹ*��N�%�|���#���X��FrmL��Ί�L���a�W�r"��6����{~���c�I����[���RQ���ʆyFb�0q�o%p��>��-������)ࠟz(�=��HW�^J3���{��[v*�g�o���]�WͿ�JT�/9�oXK<n��}$MF�G�2�LU[ �RЙ�٠�o^����ӑm�a���2=�Ț��c�+�����Ǵ��&w�����@�o����
����^���w��������O�&��o�#?�*ZI=��4뻼;ݖ�_U	8g��n='��v������5eAR�a_���rW��W�U��O���$\vn����EgL��o�MO�O3Jq��cA���9aP���w?�i��ЗF���ŏ~��)cr����<��
�^�o%���%n��?�#�g�>��#i�-BH���E���L���b�l>{<{��hy���,�|�g�֐���� �XU)s��w�/���|��,T+ë���y���	��i`��@��l�EF�8�r����!d6��1(q�e�ə���Q����ؓ+ªiU����}M�����w���i���R�?o#���C�{Շ��GY���>k��6���>���,*j�Q��YU���:q�zX�t����5��rg�����b;�\Ş�x�~���VWU�ld����y�o�^i(�h�5�������*b��:C���m�e����"ɐ�EgiOOK�t���j��ί�)ڛN|u}��{r��a�q8���J��vas{���IU&	 ~{��ޢn�`�T?:z���}�� �6H%�qӻ{�p�N�|�� j�������\[Go�ilX�䊅ѓ�C��iU?��dgT46�j���;���J� �xu��BY���Ԇ#�nl�M�4SG� g���wOJ���Ȋ��ӌ34r�^����}$����S~Y˯W���7�"�;�����̞�%��ݽ�d.��+�O>�׽y�N�+�{T%��.y���o��\��"]�F7�����vޏ߯�W�c�ry�eOX�~�7���_14\f.i����D����k1c?��IҫЛ��uq�́�+���+�>��[��=橔ͅ��r��v[��G�X���i��~���'�$w���O���1jO�el�T���5���Î|ǈ�%�k�߂Bd�z9XJ�B&�������O���*�ʕ�l��]G�;�|t}��Z�C]Lq�:�>�ﾟ�~�n��	8Ht�X��y_Ns�b����;$n�>�{��v�;��w�Y.�RܸTv�yZ�[�.�Bq^m&�����׍���JS��v��a�z�������?���3hJ��'v��~�w���ݏp�8�îY���y�#� Qe���Ѓ�ڈLw����� �F�vq|2���������{�}ɼ#���I�H���o_=���:oH1�L�ge�J#*�?i����9{�A�*J��y�E0i21�vC$�K�lڻ���_^�>�M�ΐ�կ�2X�a��W��.����ƭs������Ō��?�r������X@/��ٕ��70ٲz��j���So���4��=؞�tU!���iͶ7�C�]�o���s�*��������\9I�s-�~>��՞`�f���"�#,:?.d�ڴ;�;ϯY�F��5�`m�DՄ,E��5\L̪�A|�&�?n��D�!��E����ORa|��ԩ<�	U��÷]���@����{ܔz�9�Bgh=D�d�`ᵯ2'yZW!Շ��3
_\ ǃ���C�:%���!ظ,�� �^U]	`6�e{�u,�\���^��,f�Aґ	�諄��n��Λ�N�F��x�ۛ
�,�{˙�]�[���}c^ 	j�UF��$��UA�q��F�VQ�3�n�Gt�N�h�>Tś8OCs���GL�0Z�����̊}b���y}�|�8ڦ0P%��`�Jq1`G�|�\BQͩ����<�t�]�\��}�)M�V�I��nm�+�Sw_���5��R��5K�А���7��v�QG�N�����*C����~��s�;I��ݟ}j8��'.���i�_��-�.6{x9�i�R@�OY�)�w�hS�>�1�l"N�Ӗ)���c�H���Ɯ��cz@
�oB�e9v���l��M�0�9?��?�^�@ƕoo�l�wP�i>����#��ͯ�[���~f�e��O����E��3?5��7/3\���������Ԫ�dv�++?c�*#q��ti�K�7-�%4ǟ��[J8T$�Y)��>�sMV�k���Nӌ�T��*����@e1}k��Ц��h�S����&�9�o�ޤ�� b��x+���E�4����1�m�R[��y�EuXM]۹������E r�c��qy���j�|A[{�I�L��z��H�+�nUɰAtNrǬ�u2ڸ�T�+���������*�
.+�c�-ժ����=� �|j�������߅�Ү�F��1t��N��t5nvj%�H�b�(a�0[g�Jp����ޓxfN�N�K�[�ZU?Ik@����\�]"��V��9h�ɯع�ÂI�J���^^6�L��Xt
�&�9��(�M�V������%�{(�I�F����4��Քj���|�;*�>���5:��\:��T�"���ep�E,ެ�B�8�Q^�e�p��^�ȴ.�<|��6<B��9�x�z�-R2��S
���������g�8�fc�yxve�M6�.��S�g#����|?_ܛ��s�۰+�����;��Q9�Kg�N��R���N�Ū�r�� ����'��ܣ��4۲��G6ˤ/�S�������W댶i�ܱZi�;���#�	"9�Q�Q��}��������$w����T#�^}�t���+>Go���:��C��Ԥ6We�OL��|�}q�}�u�
,*��)���ߚ���c��}!��K�h�ߒ�����b�$��z.~x�T-�����y�K��u�^}B�E�g�'MX��6IU�Wu�L'����v�l����z�o�G���v�H�e�xpH$�1�[ީ@+t	�=t4x��So ��*:@aǞ�ْe��D�8�����j�/��m���ÓW��[D�DC�����qU���q?�d��9̊,�K
��P�U�rV�ޚ�A~�K�A�7yW���eu��(X���'�_/�̕g�w;7�%�����u��S?՛�Px��.�BL����>��`{ﺁ�g��1��~�ۙv� {�W_�������n�����S�y���ɇ���M���ت+��JQw�lw���hM��T�7��F+t���~���g���^���s>�i���T����I����9�\��8`�d\S���o����OR�]83�fqY�D��ϧQ����Ï$���|�{���?µ�}�^�Y�����Y�oD3���O��#`����Y�EE����M��c����g/f����OÖ-�)�V�}��Q)��?�J�f~�K�����ې������h���*�B-�Jl���0l��.?�k�� ғ1�1��=�6�ݶ���b+��`Kc)��D�ԤZ�V�r�w��m����yG�y��$^i<*�Kq��>˘��%�7�ec�a�$�����̣�}.���N�P'o�F��g���My�T�b��r����f���gD���T�O:t�S�z���1ѤD������ �^q����j><��B��
w���n�9���z�{C�u�z���9�5ڣ}���*��S�&m\�7�t�q	���/צ�39�V�v�^�E]9(UVż�S��7&ɧ@����<Œ�@�g��om��c-�'��1��i�T)�ӈ�E�z��l��	1*��*z6��M��_����6�Han��=ڢ@�@����̶MP���
}29!G!���H!h�l�F�I��Ѝ��q�7
z���5R�3T�Va^IG*�%S~zb��A� Q���!k����"�qY�AhL�����CMrpj��b�t#��;̜O=���uTclp��T������\RN�?1z'z��Ջd�=B܍^��M�묹�D�p�������er[-^�ÿ���#%�t:�\ڋ�՜��D�Z%�GeI��)ɢ�3-j��6��8�a�&k�2��E�d��^X-�a�@�ۭ��2��Xc˷ny��;�)��B�YCO�&������F���M�<<^�� u��j�٫@ H�~��_~����LO�1�Q�g1���۴;?M>��a�σU�ƞ�R����k�g��m��I8�|y`���"����S��-��*�)G=	��@��֯U�������8<9q�!z�۴�>��FqH2�H�R>=̛k~ظ�z�Xn����8U��u*�?�W����+�q˟��;�
���A�XUh��+�~�/BJf#�̍��:����*[n��n>;B��HU� �r5�!o���T��RV}}��u�;�'�2y_>�o!�Vs")'�v51���>��uU�����MV'�E��O��W<R,ܜIf��DJЗ������UeU�)�3��TV�]�T���O�6]>f�v���^q�����rf������bj1�f.)��`��EG�E�æ��m��/�X;�9�Γ���zt.����3N8k��s���S�z�::����G^��(��<�ϋ��V"A��Ѝ=�덳~B����~��&:u�6t����O\q�u[*�G��{�"ވ
@Dl�œx�#O��%��Eei ���-�7\�.�M.��%O��J���ʿ��t�V�V�K�[�w��Ӹ���,|\OҸ�L�:�2̅�}6g��S��O��S�ō��7}��1�
q���eEs��G���6�zRSY\4w�˹��8�2���b��(�=��|�@�sm���d͉�t���5[�vO����P�̑6U'?��sKךqY��V���[f�t�a���#���t��s�!�n�cb�v<2����i��2%���u��*��h��O��<��N�o/���_��H:��0|,��̩���%9��с��|H�%Q�Y������|i~��j���UE���.���,;N���)�m��`h6HQ�3�\�L�����UL��&�1b*�uu��L |��A�W�um�)�(�$�J�1pb����2�޻�b����=m0��jn�2�kˁ�&��M'�ql�k5?b�\�>$#��-M��*��ˆ\�:�ӹ��D~{}�[�H;S�s=�-[�r�}��RzdVZ��FW�L��d6�n�WV�>؄�6��E�L�ͺ�? ��UӃ�(a��b����pZw0 �T��x����(����-�]����+b�8ݣ�X�>6��mZ��q�Z8��!]H�J���қ�Z�r�sG/����N�k&���ƞ���� ׎j�ȓ�Ӻ���q�W�Ga���y��A��nɝZ����t�ݨ�ē��&lD��K_���$���s6�|1��O���}[AvK/��'ԌBc1�_f� |�iK�f��2�*t��n���	�r�R�@Ss��G�ȁ~�c���J�%�?E��\��;���*װ�Ko�~���ꍉ�R<e����n:TI�,�p�e$�%H\^YsK��,������s	y��K���m�G�v����qo"%-TaŞv��4�g����X^�Q���d���AG�0q��BF?���'
QWqZ��T���zf� B�B�	���7�T����'�1�3n��?x%���ܭY���V�	��{����7�����"��s$~�=H��zf���7�p��j�׸s9���|<�K �W��66T�M��U�w�=��H��(��6�jUn1���y��t?��9`7o%,����t�Ь��-*��&V����y�C�IwR4rA�����V�����7�_�2G��p]��	Ѯ*_k5@�j��y��?_}���9Xw�8f�,��BƜa�}R���r<�?p?\�K����?v����P�p�_p_A��jv����r�%��N�e����A��t�Z��oC�߸LB�/�#͢�1,Lu��8��5�B�$̤O(<���c+ӫb3��ю��)�!v~[�j�W�Sλ�'
�tKM�i�52�ҎX��P�������ʠ���=���9vE���l�YK��L%�b��W���ܲ�^��`�y��8 C��U*�p{����ǽ]�T>&�kX��w9���?����������|ס��m�#dTn�П��w7�W�ނ��B������Hq�B�t��cR���u����c3�ku �}VZ�5��:�¸���nb.��B2Z԰2�S��ZϾ"��k��
�������?���%������Z�HB��բ���J��uzx���Y�O�� ��kf~��>�;�U<�<���[��^FZ���P�J�� S�;��K!�9iUsxد����iE�fڕ����.�B
�w��Y|Õ�ڇ4'������?��~������ Q@��B�Krs0�E�g�@��䋉�R��:�b(K���:!M�*�x����,@��=��FMT���
#�/�6��X���a��7qF�)2@��<��oH]�$awL�6&gz�:0{���F���J���^�ZGޞ^�� <N;�ٞ��.���ٹ.G���%���E����܆�  ����$/R-�IvP����^�N�̡�0Gv�h�p�Tpꏣ)!�3�}�$�.L�0Mͣ�ˊ؜ߚv�Lf^����.3���e�\K�ⓡO��o�8�����\42(l����옦]P�r8s�!�R����� �>���˻w�z�]�/�v��ǎ���?���E�[D	 ��l 63�Wy@�ЫL{xy�����;m&��Sm�^�j�Ͻw���7��(�Tv��Y
Ƣ%��m֨;��ٳ��\��+��N�
�P�!�48<A�P������8d��T���z� �5�"�oL���}�6����^�jL�^$aꙵ=�Tݽċ��x73<�v�Xrjo�)��*"��m�_i���>�*1�zF��'zN�O�S�&������u�~��_h�/���HzN�9���#3����7_ioC����9'��D7#0��a��n_je;�p^�N`/�c%����=����@�IN@��o�A�e��������2#�v����{��j~'v������N��
�����&Upٮe��j�k�c�&�#�a'zy��J����z��US`sRӾx�<=P�|.�aT�\�����?�ez�yw[&���0
&��ʕ3wqް���2�'�X�s�,_�i6��� �cދ��� ��ޱ�H8�i�ܢJ��拜>����]:�8�my<� R���:�:�v ��7�K�f�R��2��f٦�/N�&7'U��]�9��1䛀b�И�d�k��f-b2S�;Fi�g�谀��r�L�z��������I��C�n�Q崁{��9&���-�E��M��B��r�.M3T���O������½Sm��U;U>�5��9��e�"}���iM�
�����K5&e����Q�)�*Dd��D�U�6�&V�Z�I�IN*�.PL����Ĳ9'6L��'�利=� ����:ʙQ=;0�M�+�ϰ�Zɺʨd��Cƒ���1�� ���	Ӣu�S�@9�,d[9  �<�:� ��w�2�NlX&6Ӡ���&�8I�D���,>�� ٪�n�!Tfi�%9�Q���p��͖-
0ܵD�%(�˲l��Jq�"!Bh��+�N#0�}oY!�a�� ���l���Y�MR%VXUJDd.�jg�R��A��G$sQ*p]�3�`q� YG�ܿ^�WNXM�ޣ��@�fa6N)�"�aޛ����k��Z`�k�y���Yr���(�7%c�w�Y�Ҁ�d�L�����88in�wY��z�!�<м��!��\oS1�uG0�gc�DX&ƨ^U���w�B �C�H�� ��)Eô;�:�	��,#�k�j�B]���eV��h�DA�	�Y��QNבR7&G��M�U�m��l/7.�v�\'�	��A��A��&�m�#v��;�~�|�gx���F�H8Ͻb���� tE�^x&�B�'N�C"�%vAJ�ƈ6D�`��9�rW���]��&�{&:��n��3%�D]��� ���R�uS�c��V��y��/h�3ܾѪ,�6y#�z��v�Â��Z5�n�,Y���o}{#�}���P���l��Gԣ�L܄+��|�x9#���y���")ζ�T���x4��Y�s�P�Ϋ+�6F�afrR7"��M�(�6٧����9)X�6�a&Jh��IR����;<�>�g�c�V�=���D)=�B$���}��!Tl�%����mt�Be9������:����T�L�$p��n�\�)�['zv[�?ä'�������7/zi�"��+"��
"HF Gru��vJpDB"8 V)�h8"V�B��3�7�*�,�pAe��e�(�D舀S��%@P�Qa�&�@�PuF�m~:4�Q.s�a>9�p���VBN-�/��1x��e�l�J��Od\'q�ܝv�sL(Y������Q�B �w��g��9#G��苴*'���9�%3k(!�4�ou3��"J�]��� �������R��Q���M��uU8#��
�a��Q�8a��"N��������PT_쑤v����읳�m�sO!��Gܱ��0��nY(�� ���P�Iĉ���L�K�<M�"�px�t�]�f�Sr(:l�c>���]�f��
&Лi�M�j��V�6@" &]A�.9� ��"rWM!I���J�ApF�!6�M��/du��ʛ&7yR��%H�$��6٩	ʥ�������!Jk�Al�i���h����J#2�Þex���=��Pվ�t�"t��������6
a�L�ktI�PkYV�i��3���`�<e3ڔ-?<Q0�[r�Z�7S�� JD�����/4�1�d'52T�x'@�����(�r�"��pS8� �tRyv9h���;,�	�pU�B�C�e��&
5��RjIc��;�hm3�`d&ʜ��1~|���䁱�s���È��ai0q^,PH���@@�p���;��kS��@� ��y9���9��^��X�XT'dl�!5ɺ��q�R�蠣lԩ��� J��w�#b�pF��=e@��2!��r�#m���O4�F�(Z���N��ee@�N�����O�=�grl����T{��9��OSқMZ��N�����9Ϥ�B,��	��Z��Q���@�"�M@3�ȕ�=S�he��T�;��Q��κ"���ކq�X��.��ʉ(�5r��X�e&S�"3@���sq��$b��X� �7)���][�� ��䈅�A�Qi:�]Iܠ��#�S$uU��.�/�v�wv@+�� �˻��S�{YXր1" ����yd��W���C_5ް70���'��'^�6���s�G�8~�����\AY Qu�Tܸ��z�n�Q+[Ӏ�f��L�Wrޛl���`���5S��6���(��A3�g䧰ɈG¤;$�7U��TriRB.q�K�.hĂA��l�+Gt� ��oN.��.y.��+�dj6� O�Z�7����&��a6!4G�*t�*��<��l�vx��bF��� ��]ݷ99��̸����	
8߰A@*�Nٌ�#�G+!+��	�yN��O��n�/�d,��
n��Q�XVj����F��≸�&τ�T���N'+�n�d%H,Xs�&r�>7��9�H[<OJ���q�l��O4�vf��"H�'��_U���P� #��O�z*��F�m�;t��� Zr��XH*
� ��_�!0�N�Ʌ0�P�(ԩ�z �ތ '�˶Bı"&���DB7DGU�Ϣ{�	�J9-yvrT�5%M��@M�(4�'F6D�vȏ�C׉��9�z:�������5P4=��a�ec��s^�.g�?��%z`��L�G'𿚂�s�!b,��Od�M��T7��,���O�F;D��:Ѯh� o�! ���Q�����,���0��$�7��R�J|�N6��!�e�YnB�%a�����Y�(�3�m�-e��S�B�[QN�.0}��N��،��Aѿ]�>L�g>
L�N��5S�!���zZ�y�U����Դ��z6�u�A�� _���'��\��\� �VX��Jc���D�9��L/6�'D� �Fa�A��;��JA�4@rh�W���=����RiΜ�:��M9��,�d��(�(�J�� ��ɁhP9�:��4��t�q�`;�"0�j"�ڬ�0Jk�Ci���Uk�A5�`��~�q��ofcm��>��(�F���Jt8�i:4FlH�Z����D\'��6�C$&s^��}�M��g$�yS�9Ѣ&� .�dM�J���`�������Y %9�3Y�L~�.V�D�Y,[��]�������:��.�5?vN[�ꗙ�.�^ۛ���h�xrMa�@ĬV�dlP$}f�I��'y�(�_>�0'zQ�!4Nq�l��LEf�у�e�).�B6@���rGD��P��l�޼8l���S��[T`�A�tF�,%Df�):�iL�WloB�������Iw�'�mOq�	�݀U?4��D\���N��#3���Ӻ�hOi.�2���,m�f���>2���D*��;䀑uޝp-	�T��ӎ��U,Vj�ȕ�,D'_�ƪs4,��@���nuM���&���e�9pP8(�	�a��<��ވ*N���U<L��r���*�H gNI��#)�3�<�a�YRo�ph��>SY�g�Db�:���2�9�$�F�� ��Z��P��>����Sa
��x/m�� �]*%Fg�j�P�N+'6ɢTP"�Ɖ�T�D�%�}�����@������I9(7%��T����(��8�%4MN��<�m�Bee���Ow��M�s�	hy仯��� �4L��1�D���bf, K�����МCp���m�$�y�L�6��<�IҪ��$gk��&�ȕ+-,Yi�9	��ׅ@쾈j(��$T�S��]\uG��)����@(��.�b�{��pX��m��c�-܍��Ei��AA��M�&7���u��j��g�����l��б;y@����c%,���{�Ԉ���sL۰�NEV�<�� ��n�!.��J���H�@�����J
�B����Q�D�x�}TM��D�lQv�n�HSPF�@M�J$��'�n��6S�K~����O��g�,���Q�|!�̤*F�m���In\���T��:��$Hܝe=��U\��豯1��6v�:����j� �)�
i�h��.�g~̕��	��A�w �i��*,����>�M�`9�G4-��nFQ1�9��*��SE��`l���NyD�z�\3%�ީ��f��(�ߴTu7:�s��j�d�^{�g?F"Q�B2���tD�M1(]��	S&�L��VE�*� �bT�D�#�� �T�c�	��o`��Su3�����]3<���Tvȼ���T�uG�!do)��6eʠ�o���L�Ú:�Л[z�k�"ж�5��O�Q~����3X�\w�U_�H�m�A�����S�$AQ!DuwЋP8B��%��ܠ�+	$�-��Q�Fh�.�i3uq�<Eb "{���Bn�ʂ2RuRK>�U7ި��ꍣr����I�d��|E�ܜ[��</�YpG3̡���%xs�L�v-�����	��4�{6ZM�A�t[�gܛPk�c\��������!BN�J*��A65N�l��.�)Vk�:��%GP׳%*S�nH���ޜ7,;� &�H�!��d�6z����Xz����������d,%���V�U�X���j�F�d��FA�	L0ڃ� "��pӪl/�T�a�k��M����wDG�I�7vzw��C��md2���F�V? <Qwfk4�	�	��p��"S�䎊�ܯk���"��4M8�B�;�_�bS<�,��u��(��܂�g��oMDn	����.�Wtw�i�4):�X\ki��vPP2�!E��sX��<��d�t͠ �3���fA��Rt��#�r��;��e�q1��<���Nkl" -ݙW���)�z�Q!T>�E�<U�H���z7�P$uXI�L!tuM
�䆫��e� �H�H+"#T�B$ ��w&�X��L�  DB!���	Lv޿�m��
�$�O�����6i����6�rX�m)�A9d�]�3��M���!07���;ѩ��l�J�5ŗ�t��7v�N�U�,�6�;0����Ifz�ej�VP�kt&sD�d�?
p��G�C�9�(�M�8BVy�:�	 ��q2�IP�B4!|�(%OJ#¨��
�{)@��a��ϊ��3ui�Lx[�e9�(�a��٦�L��	��EJ�W��Q� �"!?��U����9�TU�v�*g+(�e4Y�M�S�(��R��6�.�%0���_��nPJ �Ѻ2"5N�ha���
H��:�,����@�@qM��0=�# T� (D� E��~�`�h��u[E��Lw����`'1W�o�wE�Jc��#u��=���AX<P;�(��)�N���TsG�4�����m�V{K��j�BaStCYMj��䎉�.��|��@�Od���rq�%b�$;b��7N��kvs����RFt����T26�3M�qO�p^ckB$��T&>�Q�^�YRpl�B�:{�p:���ܻ���$�Q�P��%종�Y�&�q˂�I����e��)��--<��HN�y�U@mS�Y��
ς�ӈ"bN���
7Х�P�.!�[��4,W�F�Ʌu	�TL��!ʘ쐬�j��'T.��M�k>��+���胐u�XZ.��ܽ���K�F�����a��
e�p����(X5�b:�0�����{ųU��t�!U��e�u�Ā;�w��6��涷?h�F#}�z7�)��N�ͫ�rĶ����8��'�{��<���2�6��х<�kI��6�d�ܬ�9,�2����1װ�L ��;�r_Ü���,S�a+,�����C�j3�(#>��M��i�� �ٍ ��T�2���
ś��.7M�ȑd.ܖ�N������T���k8�c��ߎy����
��B�8*d���7N���� �yMd�����ʩ�5�EJt��7ꋉ1�8����D���� �#U����F`ꈵ��U�#�� �7�sMM$L�����jA˰��x|�-܌���H��S�
����J-�3�l�@J��.U�ɰd�]�m��I�2S���T�d+.���N]J��
u_V���C�o��Xf�r>�D)��<Ju��8&6H:�s���ƫjۚ�f+���wB�w�F*�y�1&��P'zq�(�Ȁ����Xx�<�B�(�㪎?A:�4 #����p�u�Z&���=�n�Pw��8�M�"wvbޝ��(q��HZ�D\rX�+B��H��!bD�H���D�-ώk��x�5Adu>����<�v��N����W�C}�����l�h��W�ze�pX�������6��|�C�T�:�4�B�*ޏ/�ל�GN����8Pi76U�g܅�D��2�S|\lL#(2�(%:J���7�R$?����� bT�����R�T#q�3��L,H�W��C�S<M;�@y�)�uC����"Јv '4�?w{�m�S8ç%�i�"鸋Vc�X�������x*�@1�a���T��ܝA�&l�g�i�q.�9.��c�X-�ުP.�?R�I�+��N�H94۶xJ����tf�X���N�VAr�z�����5
��'"�rM��)�Oƴ�t��>�V.TsZ*n �ʑ�PG&��c�R��^��'^�l�8]�0al,#��2�#�we�$��Y�(1;�p�� u��M���*&tB��*w5Z/i�Ay�`��4�*��㌧��7�,�H�yVӰ��QU�\�1�@\�e�EDv���XX{b�)�fL!�i�R����T ޘ0H��Q�[��9�Slz|���T�?�!��!�QB=�g@�ވ�u�vdj�	���cr5N8�t�o��*���8����&�vHoU�r2�R�|�A4"	!d�;� nS��8�Y�U�;���yx��Bꈾi٢f�ѩ@o+	m�4T�Y:NV䈈]S��@Y�L��� ��QfCM��=�F`~���V�>댏�>p��]�v:/���A�$8��5�ne4���'�h�0�eD��B"��V>tN �(����;�h�2��D�3(�@J��,:��So�Su@J�'g,�֥8(����R]��:��$r�8��}J2�@Ħ
���4�Li�A�rΨX���� �1���._.�%C�;#��@C�_�D��ȷ���.��~Zu@�;�A#���]m#����%4S]�M
��Q9(��4B:�
.S�����sC��=�(���e�����ހ��Xy($Vy=�L�N��7��%�rHZ�ʑ��c��E��c��9����V[a����ޚrP�� 
�%	�8o�"ny����Bi��T6-�T�1���r�.�~��DJ�[�EP�w�&�]�nOC³A��t�+��(�8�jքm�*�b([5 墛��(�8�ZS]=�¨�vtn��'h���x�!6�T�_�	��]������ @o�џ/�۬�8��t�K���	��_�4����Ps����ny�z�Ug�2��r!R���!T9��F�, hJs$X*����Ҡ,D"e^��a'R�u(:�����7BȂT�Np��L#%e�j@9)��4,9���e�J7W��.X�`|']it�oE���tMT�y�`�vS_/X1բ���k𒶣�!�� !�����.!�(ߪ8��l��Y4��g���6�Iq��*��A���-�Y���s�S�jSX	��ʰm=��2�b�E��(e1:�d�v�LM�Exq�s[sc��	���~*2��*BrE�Lf��X�B���B��q ҲEؑ(~j�� �[�Q$v���h�ܱ �S�4\�D�n���S����'yJ��ˉܨ<�[8�e,`� �P�@��c%�����U���24���lY�b}N�����7!"b�OwP���ۊ4[ș��z.�qS���~�9~�������8��E�L$c�5�iPx$xG5�3��L��9�p'�N-�7ށw.�h�,�!!�ʘL2J��e�5*D gDN�,���z�"T�vy�ࠌ�nN� pܰq�3�7'9���Z�o>�ѹx�}�8O�����	�X������I�'��=%�b4�4��雿��89|�I>c}�k�nK�r�x�O�;�k�r�P�x��N����r��n:�DI�����_4���ĉT��A�5�5�uM�`�x�osi��:��w~��2ܦȷ.(���E+� 7%�"�Dg��2�����XD#~�[�,SX�5G�{$�$+&�0��!<nBKSd��VQ�IN��yP�#�{lU��Z-(� 9�Ί���B��<����ZZ.�ɐ
����3�$�ᕵ��HQfn�Ue6�i�z5�N#h���� ��*� ��7;�jŜ9){��S�N"8�q`gx�mAa�۝�0��A:�u<�#�$���5h���e3�42S|�&����O�u�+�POEѽ4�%O�]���(�Q1�L�Q�⣪����Bp�����^!���E�n�����_�th�n��>�B�ru���CU#�b,��bd��m��Wad��?������M��思PT���7gs�'�sM{�WxS\����SC�rك������������:�e)��G�Nr!_Dj>�6��UłO_�4�9N�=��.&4X���w�Wlx���r��+���U�t�R��D�:��nLJ;� 5$��3F�F���0�7ܙU�IE�������\�*���_B������z$~)X�{LaX��E�kn�_�%�ܐ���K ����%6
��h<�����xjhŻ9��gx�@y9�t��!�y�f~AS��ޛ����D��4L9�������� 6��ڽ_� Z��4~L� }W�� �W���W���kX�����eQ������Z����!�G� q�� �o�]�����z����� p~��4� ̭�M��lT��ʿ��ؽM��U���/R���{���R�U"�ؾϥ��S?b&�uO2�ؽJ��*��~�vg۫�o�_g�� 2��3�/Q��ea�����i~:��~�vF<umſ����[�o����L�S��� ؽQ������z�?�+Ng�^�L� ̭�L����?���3�/���:����5�m�W���5��o�g�^�L�+Sb���\�ؽJ��~-����S=�o�l�^�O�����#��>�_{?b�
_�V���P��������n����z�9�u=����t� Aȷ��S���{���3G<O��u���{s���҃�����eI�.�	�e�
a5�*y�u�	
Q���N��uT�m8Z�Uh��숛�U�m��S�� :Y!Kmֽ?�� �F�����C� �w[_�����Wu�� �Y� h.�m� �3���Ws��� d~��m1i���z�:���_� �� �}&T�49x�~�U���C�ǡ���i�-0��6�Z��Yw�_E8�N��\ز��&�'*�ULGC�
?���� �sZ��qM����Xw?Q�<��:��r7e����S��Y>�ܛ\��*ug�'W����8��;{���2N�^�]�r.��ʡ�� U?����� a   !1"AQa#2q�BR����$3b���Cr� %��4Scs�0��&5DTd��EP����6@etu����������  ?�:��+*]$xL�'.O1ӑ���eel���p�n����w{g����@��X��;�z�t��8�B5�3�l�}7,|p
�B�mkF���A�������x��6-�����%eCs�d&e�R��pW3X�M�9u�'fZ�e\����3�;��n�_X�T�#�~�x�#fn��׌����}ZO٧U�಼D�i��(�lP��^��5\y6�;�t�&�����lf~! $,c&�m56��r1�)o���_=-��w�M1�J�'ʺ�:E�o
���c��4
TF�TX$f $q��RGs��i�)��:B�PB�ֹ��z����ng�4L�s+�K��e�������ɝ�����3��[Bt�`nrPD&9�ty�r�v�%�J�.fm��a՚�2��7*����@��X�p���Zip����ݹl	:�4��g��r�E�|�t+u��m������:J$�CD��-Ѓ�N���v��$|�����~X��n�c��Ci�or��ʉ��o���|m��ER��/�e$xg�*mm4Ƶ���R^�f#ŭ�\2�l\����>����N� �y��݇�����FW�Ы�
sx�_��ɣ�ߩ�f��%��jM�3̙���{����a��[X�0�� ��8���oh�z[ۦ%a�$��f *�X���|��mj�t����r��Z�d��V�h_^��;�4� �+!��F�o>�����'��=�g#�/̧[L�'���?���̣��	�����|W�ؖ��9a�S6���^�]���c��ч3tu�$�~���s6��A�rf�D�{]�@�{�m�?�
�SOfH�+�4�z@�]ٴ�.|0uPu��3�L�+1��k`�/�2��Mt��O���d���Ѳ��-������Ĩ�H�[�;��^�m��3US���`�/�����0#W��r�y\����J�yj������T@�����@�D\��u�����f��7E|�:�߾33�$Rj(�_�Zz���-r��㦣�?Pz�I�e�N�.�S՘�k��W�_:�qo�&sb��� 	�f�� ��Δ6��#�`X�*�Ïx������Gl�X�[���`l��H�1˫4�K2,����{�YIS�t�y�}1P�|?��ck,��Ir[�D�_ur<:���B8b��Az���3Z��7-�L~�EI+³G[�='�ȭӿ��N��/;(��kYAD����=�^���Fk�VR�S:z����$�Grt�M�.)g����#�U��&-CҀ���N�;f����ȳ �u>Ѥ#H���1�6EZn� 镆�.� �{z5=$�A5<��9�v��2\�����I>8��<:hᨗ��el��L�����g:~��{�����.`B��ۗ�x�h	��]V�Ђ��[Ruv�ck�	�7п�ʥa�ܯZ���l��Ƨ��G���5dreuk<S��j�������壬��ȤJ�i�ȋP^(�W9b�Ee�'�e0��pƏ!ZZzډ�����[�<ژ�],8ER����Y�)�=afdv6�= E� f7J��kjiY��P��,ѾSiE\��7�����d����U��$�������RJSV1��mv��H��V��<W�����Q0>����Z���M(��Q�+d���ZW1��@MU:����,;o����O�����|�=�����8XugL���S���������3�e>�w���Y��c�ر���ѣִ�.r��C1 �z�]�ʃ�ӗ�+ ��D�99�l�H�tˮ�_P+�k���Q�9h��u�ut���j�IQS�k墣��#AJ��9��͐��s�E�d
�M�4>�#�]����I��t+��S�֐��N$��I�H��kl�Fee7����I�♢���G��rZ��|��,sr������$�ǩ�o��UfU��7�u������gB3H��ؑ�$�2�,��{,q����<��#��MR9�*WB����j��e���s�q�N!K�'�ԆmW���S,F!3������������������(犲��cy�����E2x���5�/�5����;-!�|0�Q�����lFi��D��,^�1�(7��.S)��-6`=f�)L���������z�>��\�� ��54ӈ��_�{�(kK�<Aj���k�<8UT,�YjE,lṪ踷�]}�uu%��u��~��N	�u�\R����Qu��ȓ�D�e�Fok&R�+}/ah8d.���4<�_S�4����JѰͭ/HE��b��5%_����
�]�$�:s����K8[�q�i%KX䞡�������|��Z�+�y21����Vڎ��K��8��4�f����e�7Yc��� v���j	c�OО-O	+�ejz�q�����1��Q�eW��|,J�>JjU�D�i �#�%��9�T4	OJ������}p���������MQ���T��)k)(��� ����,�����
F��$T��t�c�m�ckjom��)Ȑ��Nn|mu]�܏��*h�
4?��Q��m=�k��]��n�SG=xI���s�$���"�3��.iNn����f�4SH��>�\��辰��j_�8���r*j�3�:h*��nUƠE��K�֥i���dY�Lꬱ�'R�O{!]|r��8u2�,�F���*��6R��8�}tjvU�6=bvG����1mk[(�s�_�cm理\6���B�-�#$%O2`P�Ǖ|���WX��D�i�1F���:Y�}�W������ 1��5K ��e.�{[6X�,��to�~�)Z�G`���"l39����{X�쾱+?>y*����D�@B{u5�:��X�E$�EU=!������e!5��,��K1��׆�L:���>U|ڨa�X��pa���]�q������J�ͧ�✈���":{d[m�يt��~�v�����FJ� ��X��� &�ES4u�UY��kd��.ek�+!�*�� /�m/��ن��J��=]9�:1��i|~X��#��U�޵��;�c��WE�!���ҩ)�bn� 5����dj�+h�Y���B�m
�JT��[ㄞ�����ƪl������t��J�XS-t���Q���6Gw���sm�`Ci� xxG�J� I���i���&��cY$��n���
f-zz�DϦ[�0:�</�'��2j:�]G?�0���
��LQ�B���y����xG9�� OPAP�ZF�����	G��r��@~e�Tc{�}�����И)���$��F��f��V&\�d�Erd�F�t��5��Sk;��v$��6{ٵ��hY���gF��$p#`��|�����	z��J.�讒v��0�q�i��T�L��4%H���fV���P;c��B�:Ԋ=��D�, � ݯ"5]4���҄�>aŪO��l�ٗV�ɔ���X%�k~�������F5���t��	*�=g�S�� ��i�ͽ�v���W\SQ�P��Jh�Y�����*�VT],I�9dY�Uݧ���g,�-ӛ-�<Aģ�����*ȮT7�B��|�mn/��S���?�QF'r/<�\eu�f.E�h=��S698w�����VX���m����9������i�l�4�T-g���`���P�H**��s"��\����pw���h�`j�]|`z�R�ZHX�>P��u�9�����h訠�����E�
zx�4�H�*G)gf6 `�Q4��)�Ĵ���
scg_\��D�Z9���dpHh�p%�R��r����1F/fQr���`~�q�bdSW�tp����9�o|�~�U��W�!i�s�"��C?w����{�*2�?f�h�>�klt"��i��X���(�][A�qa��������b2��R��a�	'��_{c��7Sũ?���� lz.�˛��v� 渻��v8r��0�T��}U�6gkəm�P8���Ԣ��Q�=<�j$��#�N�(fflѩ�6d�q;}!+ծ������>�=�B��{ �(�������\��?�ď�Ezjra,����
݈���\ܠD|>�YV�W2�����s��8��q�j��F�#�<�9T_����m1�&�L1/���f{�Sm�LEc��]#LrY�%�r�&Wϙ͗�3jFm:di����1`�$���9M�b��;f\�����x�g^ZK�(�� ��pzo�S�3B���U��
�q�Ib6�������!�=]:NŇ_�RL!i���I���ifǶ�YV�4ђ%�d�6�iv� .���N��H� 鵯��Da2 ��#<D[�>==��~U�����!%aEw昐��-�D��E�m������i��(��ƙ㕢 ��e�Nbڮm����6��.[������${�����r�'U�ؚ�&��&jvC>Q�$��K��#��f'���"����mC.`��w���#�9?��F�x,)i����"M��qVc������P7��d7V�I��\p>Y�����6`$m��3�rH�8GVt�̽�=���5�s+e̍q��Um�Z�a᥻�V�@$��M�ϛ*���iy`��[R��o|CR��1�$���2��l�Z�s�c��c���C%[T�b['���nm���Dv�=}q�j&��A�F�dX��|����M�Wc�E��MP�z�ʚ� �ҟ����K\N�b�͖ @_�i5�� �aP�]�_�F%6���Ι�/f��[1�����E41�}v����(R�yj^)La5��t�f�2�`�R
��REJ�%0�NFCw'%ؠ�<m}�~w���I=*o�2�F�p3�Sp	��\I,-Rʄ4JJ_Sј��^��
��ԂjI�i�i��b�����<My�&��YE�\h?VT�Z֩�Q��=F5��S���Ũ�a1J��<4�I�H�3�S��Br�k�|��F�p3e�Us��N����b��z���GN~*���@�H�NR�Z�F� ��,_S��ky����������ᤣJ���i�)�w
�)ԛD�R��:���K�D�3R5C-�]f�c_ur�UX��l="�[J�[�jjzx�����F�˝;�Q����� ��e���Y��ϸ#5�a��G�U�N��Czp�׹^x:��&��� �6�>�^)�kT��P�*�oռf���(>¢ _ո�V�����y��)ij�
�(3�;�!��PK������䨡gp���)d�K�_�zO�(�U*��O ��� �U%*ޢ�Sm�Ų��G��p_Ba��S1�]�d���7��-*Y)�"w�IijiVOe�����G�4%#�E]�ʼ��ʤ�:�\�ݹf�6+�RO�Q�H�p�,f"��9cV� ��qJxj=��Q@��i}g�l��'2��D�I�)!�ls'�J�7�Y����l=���E�X�{��i8G��̦:�~q_��i$NY���/���B����Z�9¨*��V�9�h�� �䐵�P�mh�伂>'Gi���}����H�R,}�3�~-��Y����o��l�{8|̬�Iĩ�'��nH�
IMN���v�r�d���7�3T�%n��"�3v$t�Yx8��;g�өP��fʱ����6��I�z�W�i��h�9l�Ol	2|��A
I��RV�U���8����):�*+#�����#2eb)ӂK<�k`�����T��]U�����/�$����1n�"ygӲ�m�B7Tu\�orCum����.+C$��4����WtHߙ(0��2����3���L�p���R�9�e:#[\����44R�1\�M5��dR=��� @�rBw'���A�����iޠ�c
~��б�^�� �"��v����ۂ�:�k~����"�[���`%M�ڋ����+,�6`��B*���Y6'L51
6��Z��(]b��2�*�&vԛ���pp�%5RزO86�8�T�e$��M�9��oiFIQ�
a�z�1[)[���X���iM����2�ㅽ�8<�K�kʫ�(c�l������U�.��~�+☊l���AYFSx�U�c��I�� �i.-��t����#]s�c��7E2� ���K1�G�Yl��w_��J2���m���f���!��Xf����o�X��u#$9��!�&Rؤ���rp����ʇ2�v�~��1�Hd��@_�t��6jV��R��#��:�[	r$j'L�l͎��z�_[����O�T%-�иIA�Vvb��%����5kcQ55l�~Rr �GK�;����ieG�b+�- ��XY����D���:��<����\�+?!��J��(��� �UYB�|ʮ@�А�2�� ݸ7�H�k&��Y3��e:�ř����mq��2Ri�PK=3�XD<C')c]]d���û����p{]I� �������=|�*G�����?�f�*c�]K�#>�5��,3��E�PF�_2j5Q��W��ݘ�5L�R�dK�
Kj����R|� ��WTضk��km�ma�%���'ej��f���ܴ����ܶ��I��Vix���Y X�h��(��_�zJ�:ITEԇL�KH�V�|U�����G�"j8���|CkN�������b��ş������C,S�f�si��ʌ���.
�p�1���cX�`�[*�������7�q��x8�l�ƳU�<v�x����pѸ$����MtRELXH�aK2�x���uSg �D	��Y�5�)�IL�J���^�Q�lo�l@#��T�=<�@Pĕ1�Z>[f�#�8��������H����S ����"��7�Z�QedQ������
���%-TD� ��.�����H�f��K�RF$��^uDL5�)��".0�G�.1_�+�s+ꦨ�[|��{6�a{���7�s&a �I�ӛ�E��k�����.��!�m�|.��K��뵣�4 w_<p���^�c�!<��Qrm�ǧ,�؝-�Z�QU�Wj?X���gF:0J��}��[2�I��ʪ��� ����5.�G�QY�:>l��e�t���W�U�A�'�O�G��:�F��;�����W5�Q�;� d�+�N=����<^��mM��"����c�����1�q
�h�k�Q�ͧ��(�!��WKOCTӘO-�9�K$7L��^Y
<�KI���I*^(���:�UCJ�5;ٓ��A����(��5���KIC�֦��:E�6Vs#��Ob��8�7��u��!h�f��2�]KeГ��(j�0��I��RI��}.��Θ����)�����̭o�bL�4��/�'C٠��M��(��� s9?+�v�� ���*��7&V��Dt�R*iK�1������T������S_O����t�J��(NKF��1N3ܮ�cqc�!	:�c�
���EFd���y�;��ǭ�So,qIVE0ӵІ�H2���>���`�f��~]��x|�)j����*�'����2s+j�v�UZn]T��x�<	�e.�G�Z�kؖ���˕b�Y3��,\��:��1��:��b��#�O�����ĝ�n�6����_R�i� ^������O�c��M>X�YYbN,����ˁҦz���B~��')��;O2f�\��[�r�:���\+C5�D��d�Byqc�ͧ���6��Y*U���Yb� �=L+�.���=H�6)�?�Xd������D��@�2y����#>�?��e�G��
�����frs�j|0����H�b���&�u:�[��h8�mW>�z(c�%m<r�D����dp�	V
W�ka�X�`���D[���K��
��v#�/��I�����:�{X`�e?�Q�b���|������i��G�!@���Lp�D�:xiR�:����j�FbdL��o$A����Z�����m��?٥�R���_k0�a14F�8p��+� Y�@@�X�/��x����1�����`�7�u7 �"�.!(���0J�̹V�'�u�{}Q�����VL�U24���wv��o�>��QE�3�56s��FW`���ʗU:ƿ)��|R��Gz�D\͡s{����a�E/��� ����? 1������uGE����[�{�|1O��x���!O�0�2���$��IiyyM���M}W�Q���(����Wk�,6Q�G�|4���q>Z.|��i\��FY��s�e_E��Q����F�f ��|�-O �j�L�ɗ�����C*땈'L��)��W��oZ��1u��mPѤ�]�a���bZ��Gx�pS�I4���8�A����.EQ��򭺎����v���� 1��U�Q��GR���+1�Y��EpU�]T��N��)��ِ��o:�� ̉^2�{�m�	W��Vr[&UF��	} 4��@7:�)�ǳ�o������� z���p����9���2߹�Ĩ'�Ũ��*��GUB�I�+tt̬�]N�p�����h�D���kf�d�\�@	V2�Rx��JV�x�"��,(��3�3��ap����p�YC��^M=ܠJ�ՠ�]��Oшi����~���&��'�]}M��U9'&8:s�d��{FoIj��n�*��)����U�UAT�R̧��P�5y�;s9` ]���(�z��
�y��#,E$\�u,��̺i{�b����xh韛ȥW
�e���J�@�)_}�_L�Uҹ���X灬��H�2�YJ0�V�� �+�q
8i��D��tvcS:E�WH�>�c�7�i C�E�@_�Ϸ����M_
ᔔB���I�t��f��ĹH�ePq�E�|+����Dj�+#��ED|���@ʇڠ�H��l�� ��Z�-����B�8!�7���O<�]�`e�p�?S��G7_;�|O���b��p�*��5�j � geTcy#f�YA��c�ړ��?+xXi�Ē�U�,���N�`1m� Гk��o�lqG�|J���T�OR���EG�i��	�.i 6wY�J�������䑏vfԟN�w�[�\[����2���q�ͨ6���?<�=�Z��$b��s�갵��6���*h}v�������S�"G&v͇-��-������:8f���;�1�ͮO�؞���JĹ>g��b'�ja��L�_u�K�c���d�{����b��z��
:x��F7��H�@���tgi3t�ht�=<4�\�zĺrT
�
���V;[M��[vʱC1�B�e��\�L�)�66q�T��k���fvh�EdV1��u]r��9�'�4�,����2'XR���.RF��Z۲���P���٘Xdk�%X��Z�|P�Ĩf����KÚ\����yB�]�d.��d������&p@�mX�M�[[r���� W3OIdOJ�$%�2�h�9�Fٺ|-�6êje4�U�ֽ��LfN^��mu�M�y��*^�=��<��~O�zz����l�g��r1����Ŏ�|V�-M,5��RI#E�����������6{ov��p���-g�>JW�ExR�P1IK�n�ާy�X�|���qeJ�U�W�������'��=�/v'�-�,�U�V=K���o-�>��v�Q� ��JH�=��O���#���>*�-x<�D�i�g��z�!}�yr�/{��߉z=[,u���s�$�Ȳ��mA1��_�م�u�T���I�INX�;�lN\�c"���K\��8тI��*b����2��6`����<M�êj)�%���z"�T��1���u{_0V9�c�PE�7��\RU���`��*@��m��s�`qhy�4d�8 �<�Ɗ&N�9���$���=[f��i�61�:Y�I��C��S�f�m��D��ȉ�V~X�F	�u
M�-���]M|���
9�V���#R�ܗ��C�cKĺmˍ�S6��a%��9��N؏�xw��S�Ҭ0�'P�e�\�UL���*w����qe�)+�Fs�Nf5.mc�m�Û�������7 ������T��i�GI�z�y���٥d�Y4
������ȵ�4��ݪCo�}�^�\E-.h�a�4hR֔؛�?h�Û�J��h��Q!*w��o���P���0Ư%\1�*)?�7�V�K�2��D]q���T��P��x�F�o�9L�� ��&�Z���,P#f�ݳ�*�1-�Eح�|b%���^\��@�$n7Ice�.���U��"�O*<3f�v�������Z�hEd4)Xԕ0d,^>jd!�2DC�P�H���h�<�q5SV+��Ҽ4�#B��!>��^���,�^�*Zfs�0�<p����^׿k��q9ં��̔�ґM�1�˪X�}��|�m�ZI��8�]=��%D�3��ു��������ki���y���)��0����#9K7]1 ��	�>������z?�ᒆ[�M�T&A�QFx�.��\�/���p�1��*`�4O�8yT�	b�_<J��8(3�F�^��S"uUs=����v>8��,/H�KS1s�Næ����ipUM��_��;����08��Q���/�asKrB��2ǫ>Q��B{��$'��;F�w*m���b�1Kàa�݉�e�� >8���7����H`P��{�����c�Z>#U=,t2��Jc�'��,�5�$9C�{�\q.$�X���F7s�,%�Y�п`����� ,W�<��E��-��j�4��e'�]OL�����9��Q!�F	�3#tȶν��o�6�X���"����lϙ��G�Io��7���4F��s��m{{B���B�p����W4�l��[��;��L<��42(�eǅ�؋�;�#�2~?R�-K ��d��9�r�z8���D�@���m��u9�w7���泆Sp�5~I!�ja��y#{)��>r_�/lت� f8�SH����AJ��f��xy��̪��ca�Lt��p��J�r�j�㥖e�U\��d��H��sk��_�Qd���;�G�=)���.#K��xq��B��2Ʊ��9��?4+������b�pX�M���i��M���#�r����hⓐ�n�,1�	b��k�Oȡ�Z�|���ׂ^X�%�*�M<F����Aâ���W��hݢx�A�M�c�U6u�¯�P矊�QT*�e�T����vE�A��5�!���i�x�<��_���6=B���d��7*˪������9�� �I��ce��6���GE�p�%'"���5jB�[�#e%�]K{T�Y.W(�N�z��Cf)خ\�|��o����|QS)E���VI����EWR�x��e�P�kkT*�N򩢘����D��r�/�ej	��G�����-]G�p��Q
���Cc)��+��}-�*?����=� UC�� �彷��gK��g���2��Έ�e�D�Q�_(a�V��_P� h�%t՝jπ��n�zJ��y��c~�S�����~�v$:pZ�Z�>֘�=���p1è���3��_���I�&�-�ՏDxw_Q��Ԓә�Ug�Q�����"�ͮl���#� �ƚ(�&ޱD��ӭ�GV�Q�~���.,3r�i6�%�]�b�J�'6l�+����U,J�1*ƫ�瑃��vk����,��4� }�rBԩ�����zIF�
�A���S/Ú��7���� s~��|�l���Ҧ���?�H�*>#MMUI1��⫊9c��Hae��A2�C��o�!��8}$�ҹ��#�!,%�(�#����{c�ő��*��!����H%˒�ေ��!E�=����p����ZE��iL-ɐ�f��Ym%�!b�e�&>�Q<u����<W��.�F�jUP�QG"�CQ��ZU��T�,tbp�'�P!�V��c�̢%�Oоu@|R��p�Yj��(��E4y%���<��ן@ʖ���?G�rT��*'�0V���Y�J�C��@6��K��4L��G����d�V_��`uǢV*S��t�s��F� ~8�{?ՐgS��L�?���ks������Ԏ�
��_�����lEè���㢠���I8?{�����g�`q�������C
���d�7�+u��NMt��_��=ĩ��RG<�<B���D���䠍�:Y7y6� � �s����Ģ/~�FK|�8�&߳�:YKx�#�+����=+��|/��c���8� �Y��>w_�-OO-Ks2:@��K�?�m|S'�>���~K3Z�)7���i/��a��(�����*�CUP�� J��ҡL�%���8�� X��),�Q+�	Q�c���t;yk�V��T�؎D�����ٺ�|8�2����c[�[J��\KAM(��p�+�M<��Zf�Sߒ��� c-�Xu��F=��?����S\�B��|����Be�e�2���C����%*!+��2��S�s����i���I�� ��@�����s�������^���J��ܴj�ϊ��^&��KD����x~�Q��D\g�U�%t7�h�G��{��H4dpG}�YxL<"��y|Q(�%%U_0��G�\�:6l��HśA���U�q�P��2b�PV����q�|2�.D�������v�S� 
�rϩf7���vξ8�� Ό��1	d��(5�����,���IyZ:�	q�����m�%�Y �&�A��yb.����TPL�EOYQ%FG�]��we����`���E���Q�5 �?�m�Sá�H멫^�������?25�����fS��L��j:!Y*�}RHb-xL�]jaъHУ���g/+�Ũ��v4��sn���q�ֿQW�k�7Zt�aS<�z��zN( �G>�ˏ�G%��bm�}$􊩟��>)@�,99g�M<�#}�P�ƪ�g2�\MJҵHZ^�-C3䪦��8�iZ�ɰ������qG��ڭ'���X9sI7\̧/T{�e7 �R��/@PY������k�xG�J.3X��J՚���4�*Ȑ���wt[�+�r�����Ex�A'(�!�k!_}D��ѫ6�� ��0��8 ����Zʊɞ�Ȏ7c�:�
��;�c�<V+$N
�=p4eM�>��c�`T��e�Js����A�<��oz��m��1�jE����l�5*o�k��'���IO*�"��ȁzo�k����c���������$q# �z6���M��x�Ly�ʊ�ϰ&7IC�W[;.���\2
���eF�V~�I#̌�Ĳ��m���0+�+פ �7��j�[�=6�/���Ҽ�J�o��k}-�K$�{����!,�s�6� �6�����7`�ڂ
�qko�+����E5D�|��䥞��A�m�\��A�ϧ��燅�0�ص��sI��\������4h��"�f�d��09�f�w��Fb[L����"��S����n�,<�`��b�u*ڇ�~��c��)��o��dT��:��j�S��+�i�<��,4�A,��[�G�	�rr���$P��BxsG �-%��E���+)�mlW�G�ֿ����秙L}V̤E-IЀvk�oF��� P
�9`of�}mq�a>��.7� R�+x���O/5)ii����
���#��-srnp�AS/F$���
h���>Q2�q��0�u�N��r�����@���ä<f�Ay^�Fm�MP�M���	�$W�?HxjҔ�\���{��b��t┈u:�TǪ�[1G�=s�9���]�� ��1 ��� �{�8�qj�Jհ��N�*9<�e��m ʄ��	�N=0��9s�j@Wݲ�㸿��ka�?Jxsd�h�1���Q��}˕�1C[�j��Rd�:�H슬���4=��٬A���M֒�5�UV��)��	��8�:��3��������Ǥ����q>2QQ+�5�gVȡĉ�R3YK�~��� ��W6��X�v^���QB)�Y)�=ZOqW+xs'�&�;�6L�k��,���^�RL`Q�-��� km� ��m/��KGSP_�Фld�2�|�D�.S;@�(�c҉r��t����h�ΜF����#�qs�V<�H������ #��0�qf���)�ѥ�{�d��7�����<�N3G�K_D]��M����f+Uh�<�u�
�����3@��>��"f���6n�k�5�%-��� h�#	��W�qulþ]v�=�_�T�;<{~�N�VI(�*� w+�b�Zx��.o��Ois���.���zJ��i�l�:+I$M�U{4E�ʶ��+�� ����S��UW�N�լyi�g�l��"�WC�	 +�x��-L�Vt�`�ξ��#e�zpZ�"Dy��C��0f��V�JjSL�T��Q��a H�ӚC�P��:�85L���X�z(r�)�z_U����~cvc+j���V��W���Oqm!�����ƞ���GV"ڿ:�Z��x�2�ɖ��#N����X%a}[�� I��+�*Jw��T�q9dn*Bg�C��9�gߺ\*��_��q�?ڠ��#��1�0+��MT@���H�@�q�������<���&l����!�r0�l�����=,��^�N-����+���KC�Q��{c��S(�R#����C�p������p�bۓS���w��EU�.ҋ6i*z����2�������^/G��?��K5�<���4|�:�Uq���#B��PIFޭ��R�����:�������J�a��i��^�[f��1���������F�Y�z�?��(y*٠�97�S��;>]���g�l�H��Q�L���\�	IG�E�	@�$hO��J�t�>�7͚�(�Bwǥ�����OySɣ/���|p�-���σ�h�aI��٬���!6`Y�@�۪�8�<A׆Dԭ����5����E��>f��ks��P#�˂����Qu~���;���'s�\�8RcF�T�J�Ȳ0}�t�S�%�4��1>�E�gS�$0�am����2��g#Hs�r�G%P}E��-��C]�j'��{'/5%Ub�$Ϙf �����],s&+8Ȧ�b��L�	u�?)�����,��v$rx�*L�AԱ�ax�e��� 	�Sm���Fi��I&���M��#C�[[}F�H$�i�����f�!y���m��GLz����`rN��)c!y�w�ݐ��ɓ��w�oV��k���<c�UO�Z�U����\�Xl� 7թf��<w��s���PeGue��{w;c�B���G�A�MX�z�~�/�k����=��X^%Ÿm^HeI�}xA(W��ylTH�G.b�E��ZO�)��D)ǣ�='�qtl�����]�G3'� a�^^�xuM�6��̐�����5��[�q�U"�����k�c���iK�UW<<�3"�������� ��$��H��:
iZ5l��/b���F^�bRH��&�`lF�c.��WB�Z�c�zT��sRFME,����塨�syQ���Y�	b22�Fm8K�X�|$� �Q
��ǘ��k��+:K<��ݍ�~8�.�߁�D˿���L��S#��/�(�x�3�bq��Nl�]n2��ܔ�et�����,sR�[��Yz������pde.,�*����S�{����k�K[NZ��F II���K���c.�f�~�n�J�?�&��/`��~!�2��K.kl؎8�s)�b��l�.�!Kls�� ����� ����:�y(i�U�g���=;�q+̧�d�)�=����Y��}u��-d;i <{��E�����l�L�hzCoo/��k5�eE�l˪�����n�7�ت��<qO\К�caʔ�ư�r����˶��z�'ի#kJ��ʢ��kuc~�1Le�����Oo���]�����ǵǣu�L��^#����g&a��6�@�X��4RA��0%=;�Yf����,z["YdT]���}�67������ ��q�h�DT�
� ���h��K�.����A��J��KqJ�?1�55q_|�Q�����tg}�j��osl/�_��^<��?Y<΁a��F,��h�n�5츒�h�I��B/bG}=���2�34o�� �<t�?�X�bܹ��$#��qz�J���|������	:������Աǥ�����QR�c�I�_U	?x85KC�_Z���/������43�z�N5맑���t��?J��^�,&d-����?n"n)?���Dke�������,Q3�[-�q�&�����I2���2:<L��R�� �G8]D�_�5ÈS�Q��4R�f�Ԝ�3eR�2�e7N�Z)F���2��ΌȲ�,�{=�!�} ��H������Ȧ��Xv=��K�]&<��2ϖ�W`��o��#�J8����<��o�L�c{2�85s�˫1ċ$SH��<���r-���6k�?��u�JZ8��LT��D�_W�&E9L�0��5�7�r����j����+�QMU�hퟤ;ٿx2a��ߥގ@#�ꢆ�/�1w[���u3ils�.?�|"׶��)���������j^;V
rh��Y��l�B<��)��%�?��#~�� ��x�:�5tg,�I|��U�l�X���Zj����4�	�bb#%���,�I�Co"��%��[Px{�f�h�bI��� }�e�\�48�UP�ѵ}�� ���H��CB�Q�
Ŏ8�*Y����m�p�m5ͧ��8���Y_I�h�,�T�N�X#�I�fʊ���:���U�SEPNu��*�r7a��8�q>�b��BD�t�1�C�� Iaosa`t��� Pq�W>cëL{����;c�է���'���y��YVIs���nqQSP̵<:��jtE�̴�m�C����w��5�Hx�;u��P�!ʽZ�7������WO�T�X��YK�O��!khX�8��<?�*^�� 6����L˚#��g����6�HČ8W�@}��Y؂M��Cm|�%�U��b�ե,��BF��_��U'�C�qI�*(楚Jg��W�c���&ev�������a)��h$���J�y���L_����k[�f�n����d���Kxi�|RPM#�>���"D�8QN�	��\*�M1SL�u$�/L-���q�������ck��o���C���@M$0��J�}��n�m�V�u�Ds���u�2!�����b1�x�����$4�T�ai�F�L��r�e6��k���,L0���`@��r�G]sf�G���4|�_I+���R���N#Eɝ��*?�{��
I�,�ᛤZ�y�.=�c���ia#k�:�s[6��ط�)�ja�`�A�� 7�4K+<1�$BH�A�6����O�A���c�]66
4Q�� ����R����ˏ+��fӵ�~'X��$j=\-�����!��S�M@J�Ӻ�-,�&�lF�U+�w���gC$K#KL��@�e 5���_y���Q��[̀1q���I`/v~	�WR,E�����Z��i=��=�IP�����z�HtMYn��O���J�Ⴁ��"��2�Gw�ֶ\TNM�R$�E�������������[�<MK,��鳲{N��#� %7�G.gOgU��������@_�q4��ă����������uc��C�i8��2-�1�E43�#7-/"뙙�\��u��>���g��_ִq7�p���4����\�8f�u$1чZ�ؗZZ�Fj**�G�}b��Q{���;�Nm��J�������M9V��6x�d�Y�k��#髸	%,$�f��6�|�⦳љdX�Y�9�0̣�I������
���_��'�*X�
qh�f(����P�c��=!�U+WG[Yϧ�E*��E��9���Όqg��થ���𡨞XJ5C\d��2Y�3+=�3����xD����MD�9�˻(m���툅O�f�R����iV��Lϔ|�l^z�F�l~͹����N������^��pZh�ܢ�QƯ�s�9�u��01�T�b.���-���}'XRa��������$�Zh������0N\�T����N�mz���|K���PV �e��fK���ݑ.�t`A���8��߯e���t��0�i s,�!�Qe'/�A��$�R�Ѩ*VD��L�2��_���p�,o��5EB�9=�2 �Y���'+�il�+���Z:y}L��$`�Ѵ��7ao�⾾���/����Y�h�8�*0ܜ��y��$}E�g�����^.���z��p������.h�e��9gl݇��O�'��iT����DS}�:N��FV �0D���A��X�����G����?W����[����"�Y@$�5#>�'�ʧ-�e���Ԛ��lu<��2c��X��L�GOP �WIƥJj>%B:���	���Edi��B�b��� �N)�}+r3�2<�3X����k�'�Җig�g ��k��bA77>S'�9�Y�{\���H>6���E>�|�%!~���z�#��>��x,.e̲GSF��e� �s|t�8_�|V.#P�bJ�U���q����S�yVoe�E�8��<;�p��R��
�囧s����N)�Ӌ��TVH�d�5�<�2�|G�Z��Z�M_�8|0���uk匳���t:�}�U7�+_�sNu���9i{�ok`�x�{�)<�ӗo�Ⴭ���`��=;�!������km��盉S�*��"H�W��J�"7nk�n��{('�����'��c���)`9YU���H�0�{� �܇n�s��sI ���s�;��6�ga��e�l��^���l����.�� �>xl�Ë��KGu�p�2;��J�!K?+4Jz~���x�~c|K��&������T3$B2W5��$j�̥̤��7🁰?��Hx�?���"i�j�`�s�Wf\�b
r+6^�Eo�~�Up�Z3BRN|����e7�[(+r,oܯ�������QU2HYՂ��t�2ϑ��c+Yd]Ɲ�ƾ���5��)@� )� � D�����dc�+����Ⱥ�lN*8�h�j�%0I���T͑@�76)}�x}-���6)�(h�����΃�$�@\ߓ� E�*1NX��Kg�bN\�ak+�䧊9.&�����p��6!�o����2��bE1��R����+��xbF�7�������c�����Ź��o�����]�?f?{1� ��¢p<9��͹�c�qp��I7��'�R��+�6��΍2Į�2�[�n�K���Ѳ�~euQ�X�.nh@�7S�Y����L��_�ý���xә?�H�6l��wʢ�e�w�eV��z���H���*����*�	�7����asp� C�j�,�۬F����AQ��n���V�v���J�N��I�x<�S��P��S^��d�7-����|���\5��:j��FHa@f��}l����r�#�����.���a�1���-����!����]a��D�3���ZwuSnĭ����\�����(�*%�c���3�/�fe�kk{ckyb�u#b/p|t�p^��1���/.8�FEi��P�-�����L��
�i��,1-�u�T:)����_e��;�`Dxl-�[K}`$(B���8-� f
O%j�96�PZK��{y�Z*%���-*�|t<#���94u���Ӗ�R�o���Y�-<�$S�#�4N2�R��7S�tp���E���Ǽ� o����q��%��p,�s�č2Ŭ��Ȳ͖��k��.gc��qᆋ���� ��z�J#�f�
9V6�M�8����zM���V�����{��}q�˷�^7wF�S:��T��bxr��\��� b9nO�i'�%o㒐�;��a�㧣�5 �tuH)���s2Lcx��#\z��&��F��YB޳(�nj,3BA9�~lquf�Po��:���[���/�� ,\K*� ���s%�[�H�����g��,Ϳۂ�]V[�s���|��c޸'㘶�9��ϗ=���ƕ�aN��D����m�Ү��� ��?�������rA�*+Ҿ[�����AiQ���ܭ� �e��q�U¦4<�t��aZE|鐗L�Y3:��a0�Cl���g���s��(LS�KPY�=f	{$pH�"#��8}u-,��5U#G�h@�Ȋ*�9]j{���٢i'�CrVK��9T��8�mE�M��xLz=���R�9l,O�25���)�#��Ѵ�<�M$i:'Y�f:��Sc�1�W��E/���U�G<�eyQ3
��e�[�1����%-b���c�"��h��V=BBt��"�	�aw�)���� �J���nc�O��,M�}~� ?�V�W�~i=n@�t��h�9/wS(��}ˋ�?��� G�?E?�<5"�X���X&�Xd�X�]c�H�4c����s�"�k�����ÏJ�bt̆����qǸ]�����rj ��nڜ�/,��*H��o�~!Uʊ������9t�9��T��'-��p�GMQ���<ՂKIv�D1<y\n����>ǫ!�Y+8r�T!��,N@�wL�r}潀đ�������X㑤�	��I
�eUuIJ�X����K�'V����I��J/"	
�X�^6ka��x׉K�����Fi�ʎPT��.H�3{1WEƖ��w8�����eZj�)�$��ɑ��9��4n��z�����ü����o��fr�4�I����TI����8��ʑ��#��y~�!)b�O�ݣ^ļ�ᯨ����*(�Hᗅ�IMMP���jjc&'�srI-����)e$��N¾�,��$2s�UpC+r�#�o��Dу��8��	wAY%=�Nk<QU:�E��V�	��(�U����2ΆNZe���BI%�X�� ���p�"��"��E�.~�mYN%u
sΚ]Fay���@��5����
�C��n�P�a����a�SB�#~7�X���&�2o��m�����!��)i�4���[��g6E��L���R��8 ��L($����ѹJ`1|�K�9�7�|����o=(�&֩1��%�b�u|������X��4��n�s2�n��NMߘNU
6�*8�/M7*�N!MX�$�3@���O-�st�:�_F=8�2�C�%|�ke�s-=L�,��\J#u�n���9��} ���~��Ʃ�4����ݬ��sf�])���R�;D_��:t�$�4h�5���Cm��Q�<o������)�uk0ua,}&ٗ���x��(kf�&�{0�(�؀@;��bE�� �V�2抪�����9�7���#mp��(�z~t�"��%��+*y@��!�&�u�z�dOi��<�f˟�KNL�S�دK4�m���H�ψ�!>$��)j��z�/4�v�5�����[mb;� \p�.�+Ө�o���8�5Ӄk]KG'O�v�b�ў"c/PR��)'���+E`,�s�OVgp�$��D�EKO4��@���:�Ff*y��.��E���p�~��k��5<�)αG�)��V0�٬�����<S���<-W$���2^��T�ߝ!I	yI�a�1�(#�%,�8ѿ���m��*)�O٪�j�>Ԅ*�ʐ\!�����%\�\����������.H���%�.�t��l������G��W=}7�� 2C;2#8�%1U�ֿ%�Ą@�+�S&H�袁M�U]�%���^���/�������r�7Ԟ���]���'��S6T���'͹̅e;0=:\q^#����յ�C��Z�L�
s!��P�v��V.�II�~!h�Y��*K3%�&�������������8}?��L��I ����R����k�����ꊎ.�Ʈn+Uh��F��d�oN��d�]���f����������� JfX������ ���/F�)�T�-5;Z����2K���5��pȞ�1d:��F����?��$���B�!���D>���й�;�:�r@ľ��?D�z�#I!z�U#�Gs���@�tQ�ׯ�p�;[�5eK� ��~$1E��ϟ'Q*�����YP�q:)`d�I�d[w��������e�i��x�JW؉3C�:B�Z \�s���ft>��:�tiOT��t%,�/����}�0xr���j�k�I����TȄ�շ���Ǧ4\.�����q�!j,܅�E���O"#��U�1��)cq���b���&z�yJ���M�\�s�KH�EC#?��s��� 6@ɿe������e����õ�bXǣ���Vc5:�u�c(Y-mLe��[b�n;�'��?D5H��{�6�l��,�s��̪m�gN��������N��PL��� B�@'��U�ch��WC4r�������҆���"��g��M77�%�XU�m���5��n�Vz?G�x`��7��N�� rG�L�
��$GR�;��\p� �_�q~T
u��IۇΠ&��A˕�%��hq�(���83�,�tq�r��NQ����>-L�Qt�X��>kz̒ 檖�,��g]�O��
n��%WWW�fr2�wy�!o�c�qz\ޭU�'x��R��+��B.�ʟG�Ep�rT4�qY$�Q��z� #au�t���� �Lo�56���~��*NM�<N5��<R�d��3g� "2!��QQP�z����y$���*T�H�el�:@P
 ���G=}{�<͝�gNAbl�"��؛ SSYQN��(�� ��Ik��&�R ͨ�_&� \P%�墥[^��-}oop��'��I�m�:��� ٺm����T���igS���.�k�e}E��zN%OA[ĩ_.Ig��Z�n[lq�f+��"嵎@F���Ԙ=Z)�*dZ��34��u���s%�[0��#JKYI��s �)݊�5����rҞ�9��Bn�Z8mw�gl�������̵��%�Jyfd�(��a�]�2)��#�ױǣRV��Z.�X�� dXFK.��Q����uk�S���>1�e|�$�y��:�Tث0�X��>&�Wp���g9�f�l����1]5�8o1g�2A�u�MQ�܁��b<-m=Z:�Vn%F�"���k,3�P�έҎ��]���Q7�z�D��pR���g,��.Sև}W��|j�UE+�ehԆ"��{��ƪx�����)U
X��'H䈁#��2�7�t�	��X]��m���.�Pmm�U�~(]���P�s�A0VF���c+��?�|ռ����O�j槨�V+�.#h�nc,�]�s�(��7����b~(Yc�7̓��P͔<9ϴ:b���JFl�¯����]Q�X�!v�������6�T��TRM'&�%Z����Rk4�<@����X�l��ZS{�ʌ9�k�_Kk��()3����eC�QDm� ��\�#�>XN_�ޫ�y�M=/.2b|�gVdUfl�{ȶ&�|ޒG�E]L>�4p���S�j���d)\�HL�|�%��EO���%�0IjX���J� ׽�)`��Q���$�Ϊ�]	��u�� �N�X��eo� �w�O����cѴr\��Ur짳f������?US�P�biC3M6h&I�1�9J�1ٮ��X�lpV�DBI#�	U���$uk�H�\���|M]�Gĸ���Rr�kj$zq���p��wpݰ��%��>!TE]lv�)��mT��s�NX����?�uR�$r+TD�uq�B{��.=H�t*�6+h*h��z
�*z�	ϗ��Tc���b��ګ�)��:���~��3�� �L��n�i�ؖ�.7,4���5�!檤���tit���/��a(8�g�A�(���9�/)Fs}E� 徸�� ������=,b�:���D�(vq�d F}�|:�E���5�������5$uQ9�+��c�Z���f:yaA�㟮2��jVb��u��'^,5�S#CPI�h�c�]rDa�h��I�e��Ӓ������ ^�������pjl��N#����zJ�밵�,,
~3�/�+��*���X~6o�mҷ7������@�����F^���%�B��*C��� ~�$w�� \�VJ͙Z�M��X��SL�Ŕ 4���%5j���/�|����R��{�a��������bم�/�����zZJ���Y�\�9�"-���d�1錿1�
p���pظH����D��#�����Ĝ9�����MX}eļ�vjP�x�DdŒ�J�e'c�� ����⊴Ţ�yQA��`jǦ$5�k5�Z�+��=jE���*1���3k����lRpZ:��4��36Nk�ٙ3���<�]6 ]��֊�z�d�"��=,VR7Y3�����˝Ⱦ)}�5/KUIp�Y��EY����X�(nk��o�,|�=%zR�ͬF������W x��e�GPm�^�	�A���ޢvp��OP�$Yc���\�
��j+�%i�j�y��Cw�I	gv>,N/�~����>/A����R�h`�6$>�$�;�� ጺg]G�R7�����h��p�����[@1��0Q��E�� s,*�L�(�4aP������U��Hf��5E$�� ������)�7<R��Rc9��&- h�@����J�.|�����h��lt�PŜD��F9R%~dl ԹC���>�k��yc��w<��7&�{��ߨ�4�W��&)��%\5Q��<��0�5v钚@%NLy2,�"��鸭j�4Q��(8�ʊJƷ���6�$"�Hu\-o
➦͙R�9�%|��lZI�$�[7-Tj��)(k������`�t�%٣T/�'{o|p�98�5=%2ѩ���12$+g������D'����W�YEW�姧�N�r��"nd��Vb�s�g[������ ��MMRީ.��X����uk����i��hH(̶��gV!��Ho 4�G��ER�}[4K
���@��`��.�}�݀Q ��n�{mbu�?��1�=�z\��<���� ڧ�q�9�`6��������8w9i�ue=/�:�XD�*s
��_1툦���D�,u4���E���6e��Mʹ������ �,F���^�$5r,���-ѭ�4�3UJLn���#���"��^���o�8g��)$�3<~��]b��(
����Η�O'�<>3*l�o:�>�_�a�Fv��
�H�k�d��դ�������|:|��Tq:���djs2�O*�)�^9���N�a8T��<����9J��E�OhXf*-�����Q��X�'�Af�i]E�}v��K[�g
qarI0� L��3�Әjr+��lIL8�d&OUr������ɑ�k�+��t8�.!�M,1��#]!�N˙FU21�������!ت53��/�DOU�Ԇ!M��?� ���g9��r�ⶢ��n"ޣ,1��)K�)L�e�f�b��r�w�E���i I�JyN�B���VK���� �i87�
k5TM �Լ���>^N_S1#�m�?�>�����,"B��4r�����m�l��R��񵪣����)y�$|���,����\�3-���-m��?������jhi�<�
��01�9r��(��oz��"���.3��!�Z�j�*e��4��c^����W��F� 2��l�|��]%��~cJ)%��S��C#f������S�E˝��*ɪy�eUa#�@�"l�̬v7��Ixm4+�"IRd�G��a��.{�bHOz�a���i�)HT���}��A������q�G��R�ӤqT�P�^�g��,pH�2W��{_?��b�j�=� 쿅��_LSI�+8ubTK���gv��[�#C����i��� �.ca��(d��౷�e����D��.|�?Wk��p��ĥ�-�A,���,q�v�P�B~�b1[=�$�/�&�Q�Uͨ�(�j;���7o�ًe�6ɷ����ܝ��� m���^��r�듈A_�Ϧ�4BQr�h�+�X%�c���}i}�/ �X�f��Y@��|p[�q*��� ͜� +|�>~��:Ow�w���c��P�%��"�r���ȢA��"�lN�r7����◉P�5o��)s��JT\��T6����a�2������?N���}N)D�ZTŉ*G
���Ӝ�:�j�q��Na`�Ǔ,H�X�Hh(��������j�"���9�4�\�ٲ  @m'�Eex�GΥ���u_{@ulp9��$��)j#Q�f玈�ZUND��;�0@y�7s�H�,�d�[ո�G�
�s�T����#�#��Z� ��`�w��}�kj#��+(�1N������Z�|��|����I&T{�<��h$�%���E77�+c�x���E=b
eL�*��s!L��_j<���#z��O�y�u�m��Z��-_�fO�)���T��m�o�*8/	�j��E6J�-(��z��\ǫ���Z��>%���=]sz�����1�59\��Il�r�F����T_[��TU�ȩx��>�V�6�.c�Sq_I�*�i�hA�&����R�MԲ��|��\�Sn%K��b���.�,J*�M�n�b��k����?v���ĹW2Aĩ�43g�H���� lI&�����-������>�%��Ig���+�L��,0�B"��(�]�1�0�����[sO4<E���1�Q���=��#L��a���4����4�fD��%�Fe�A[�P� �Ҷ�KD��#)!/2�&w��a�n�m����;� ^ؠ�T��.-R��{u�jȏM�D;��rΛ"�:�U��C5	�^��E=�L��%�uR��uFL�-5W67#�1�� �[ܛj0u�ا�<T4rP�LMJ�I*&og{��"�(`�ȭ���(����O�Z�(j"�Z�z"ch�P4y$^��:����y��qU�̎� H����V���ֶ�X]J��4� r��~|pv8��6���ƚ�Ā|�4#�}���� v���m��G�Z}����(���1�^֓��n�a̒�W�t� XmO�5���?��ċ��-���|g�i���e�a��v�;��g�h�Y��#�vND1���r�#Mξ-�\�M��m5 �s���jXx��L�,7X��@�J���ьyY���X�r�ıc�-����p���q
G?�6:��q|����(k�y�y�����*�\��
薐��G��P*=^��X�ʫ`�$R����t��\ܑ�Lq[��g�s#��� ��pڲ�֞�d�2�e�k�68i�Du���sp�f\3i��.�$`\0e�9Dj�XŞ)�Q�Wfe�1R*F��0��k\���\��������I�3[�`/�[	�Z����CR�)>�0x���N�!EH��T�89J ˔ 6����$���ȚI3�$еF�0�>�P�l4&��k�͔v����I#����S̢H�y��C|ʽ�M��?	�մ�n�Ri�4UPK$�Ş�C<kP��֌���$�ԣ�f��L�i:����yXض�H�O���&E���F�ʄ�*e�]�
�bX��
�xx�]�+)j)�����x�9S�#H@���������w��(L��P59ʱ�9U�d/|ō�!��<.��p����7�֝*�����N��� Sv��:�����u�9G�-3����;�W������śD<�S�Ѯu@"��a �|��E�m���u%d�'	4R�U�2K�^(ldB#G3��XgӺ�SR�>'U���V����1�����O~����ݤȨ�	�6V^��z�A��R���9N�[/������K,�p���Ӄ���������b�q̐�/�V��YM4O���9���� #Bײ���%;E�o�Q��ec4��� �o~�8?���g������P���*fg�9��H�XU"�yOHC�S�ǅW"K�<��Ou��Gke�X�ZܰA�#�*j��e��ChT��rdmu$܌Pq	}"H�z�:�ZR3dl��.{fԐ��nW��T�U�od���Հ�qڲ��,CK���r���b3E�+��6/��t`Gl�M�S��;y�b���H~��X�PSF�,�1,N��},{/Hk
�hR��Ȗ�e����OHj�{�(�ͧ�x�������j��.9�
��4�um��_��Tǔ��4KL�)���R�m��^<0h��g,�l���,��� ڛ���� Z�Py�"��mm��Π6������%�aJu��n��1{v8r="�"!2+rZPvb����2%��m���+Ҥ�����z/-d+�l�J57�lG��V=�_!b�� �rd��� 1����J�y+52���J�
���X�mtq=C�?YO�i�f����%�)�$����+�b�V�}qs���7o�潖 u��V��l%�������<�S�ԝ$^��&ڝ��6 ��lHk�ƺab����Ǯ҂��-���rdɔe���_�	Qcħ��77	R�سw� �]!4����,1kfX�d/,�qc�u%�8�A� �f�m�.exίr|�&`@m��i�S�s�,9i�m��f#7݉,��3���LXk�e��k���O���X�E-wꨦ��a"vj`}�"����[v�ؒ�GVy��~�Wfk 7��[qbn܆�~�X���"[��h�P7,�[���t���)�$�*�/����-�F�!&Ǡ���6�Y*�MF'��w�(RN`�۶BG�٫�x}��I�J���U[<��i���n�zj�H��t�V���`��*!1#rң�S��A���'�M'x�H������H���,vl�$TA�x�L2ȱ5��6�x�D����{b���Z٨Hл��VU�� "��%�r���>'�=r�Ұ���J܅��K���˨ˮkSx�l5�^�1_��
�&�[{^�eN/P�Ւ	���"� ѫ:e�+��c��k©��gIi�0e
m�(�"� �P��\K�JJ�ji��Fa&T��4q� ٺL�U�6�)]]P$�<��z� D�X����eSp��d�QS�!3z��s*B�3�ic��f%6	��f���AAu���n�"��kh���g���5��Ut�!ː8�Oh_)F��O���+$P�Gfp9�W2�8U͘�4�u7��5l��9��}�2ʑ�-���f�p�xut���KA�-�M��\��;/��J�3OĿX��*
��ek��D�I�P�EJ{����-|,�������� �ث��G�I+/6*U��&�2c�i�)mzei56B��ʔ��6�_0ЦB�Q��*�#�������#�Fz��������Z��1n�b.�!7�KP�u�|�_u?�%�Qj���{Z�l��+�u���髿7�5E�3
eb��s}�>bm�����M_ �4��z�VJ�,�K$@ك�ڶDf}����k���E�fz��6����2�!�� Qz=ţ�)(���̎`͙��:5��mf�5��\l�Iq�3Sә9AT$wk��P�2ws���:J/��h7�$���K�>jF:�ڞ�����}��+~���@��-�]�9cb��|�l+�kB������$�5��焢�\%*j��L��Fҳ��r����ˠ���f�ε:�l��	�3�l�[���6�� �궣/�Zho� p|��1 <����2�sN��s4r��b�Py����5p�§��(�e�Q@]=�����]�`~'y}^Fi��1��+��d�ўֳ�������������|f^#19��䋁�Q06�q�#�^R�J����岄u?U��P�{���s��)��?]EY�X�(Yb5�/l�MO�\�QI"fm|g��v�Yd�-J��X��DegL��l2)���3л3��_����`I�[i��6���ꌃ����(9_7,��u�� ��_��G��H�2��X��0��K���|s�������L6f��V��By�^(ͯ&�#&�w��b���9�\�eՑ�:�-��ªI0�PO2b��1 f���*4���̊Ϋ#���!Q�E�p,��lO$YM\�U��s4$e�\�p�A{~��VY�tN��2��t���\ub@-���q�Ӿ�?r5e:�S�s؏��ԕ�<+��Q]L���J�����,���UDd8U�7�[�E��E�>k��9sv��
yG��QT��r3f/{t�/����2��j04���Im{�H����x�t��?��GFH�*'���˒je������RSPR���I5=�=�hz$�D��}#V������̏3�h�E.�,�]:������Վ���P+��-�%�@��MY�^�:�%$��
ML�jYNn\S�Yn��뫌KC��g���K4y�B!��,L��%�_vU���|�������%��X�4�!�>k��#����1+�n�Q�$�,yJ��#)W��/���\5�DK-��gW��.C�\//������C�P*r_�Q���Lel,�S$���(k�'̭�|�o��>1�)�w�Q���hԣ)�t+����I�i� ̌�,�{ۖ�S�U�{����6d��f�`�o�݅�� ��5Fd��ȱ��BoN�[8[�e�mŝ VD�3&]zd�v��|s�qy8�=m��	��4����tAo<	}~Q��.*5��$�/��V��$���K��J����$h����M�L,P�(T��ʞ�Jo��S�s��o�<��%d��-h�#a�P}��t=�} �	�d=�+PJ2�_��3[���+}�_����q���
79M��}k��7WR�0�x��.�Oc�9K�#��~�� Ą%�=co}����{��+�ѹ�}j�'@�f��h�݇��~*�F�)�H4�ّp/�p4=���U�K��fN ���yU��V��7 {n+$��4���bm�2��'1�X���Se-@�dE�lЯ@�B�0����S���V��r�/e'�˷�/��-ח�,"=;�`d�� ���!�� �z�H�c�W�d�?��������N$
����2_��f�����ę��R69�|�.���Ƕ��3 �0To���}-o�Ï׵-�9�e#pn$Tj���?Uh���t������N���$��+���Cym�L��;�\�������|��M.4�}� ��âaW-G�V-iQ���Ȓ��n<襩P=�&�S�J5�Zv�K�-��̍bFFQ�H�M�s�ʸ���~�'��e� ͮ����հ<Ys,���Cl���y��j.r���8z��V�|��L~6�����:�,�Z��F=�Hܵ����$�^�$�\��! ����\h�Z�i�='�B}�i�KYIb!��v�9�2�,R����iH?����&��_[�a��kk�̍�\r��dw� �5�2Fm4�}��1�h̷T���f_feAI�s�F�򋰟��:U�&Y)�Q
��2+�U%�fb�f=hڟ�	��s�-	��*������<䋒�(;�F��H �GX3$�*US{�W�$X�\qE��	���R��J�xcXƃ<&f���bJ~߳q:y����r�e<�M.^6kn���!�D��7�:��1w��	5��I)i�fP ��%�O�T�����a�2-~�Р"�Mvx�D�a6����w�����OY�/���2-ؗc����������	�Za��8�ȗH�7f̪����Z ͂?��5�m�����ʨ'`�c���
`y�r^�9=���ǹ�FP͢]CZ͛L����ǣ��Jū���'$�`��v-�}v��|��K�[�@ya��6Vܭ��l�]��0�%[��}~��������Y]�����/ã^*�O'>2ƚ�"��p��Q��l�u7��J�*����2E��$o����̍�ݹ��:�ҩ�7T���� �tч���Q�y��ua:����V�{�LU�y���Y���3�-UP&
��}b���B+2�#<��|T���)Đe�6���@�Y�L�Q�$H�J��ʚ����/�8��~�R�����SpŏNs���%�dU�#c"��
Nb-o��, ��|�8�D�>f�="L���\J�+��h�t�&Il���F�X[TU�� �W
5��u�ozױ�ë�� /��f��Xi�EN34k� c��j*9�l�_�>��rⱔv�E�X�/'��T��J���]c�k-���k�hߋ]c�'�GHR\��sO$fK�=W6��꘣d�JR-b
zĉ!n�_n����x��k���}%������X�^*�Z�1�CZ�3o�H�Z�S��O3�� ��IM#+�0�Y��vg�[��G�$���gQFJ��$���[(�r0r�Tʙ��&P���v�Q���Ui吜�d��h�>��*÷A9[��"�D����Ypf�u�	2�X��,�����/.A�IR]��m��c��ȋr𹨫�i[k�VG���SD��5YU^ ����2�MC���r�-����N���B�ܟ�ꥊ�s`��&BW6e��-[Q�d%�v��^	b �6U#�'�^έ�I��3ȧY�����48�5l�i������X������|f��y��%C�Y���*�{N�uˮ��"�OC����^Vo{[� 
���2R��_g�3[R�����W,i���؉Z�,���9�S��r�1}2��S���ꜱ�I���f��K�a���c\�q�5�Ƞ������ +*[�BJ*�}�n{��Zj�d)�D�$z��0���a-D,��?�O!$���Q,���L���V��_�ҊeWYxIhd�l�.gekx���/�x���
J��3��Sv)w9C2:�Urs u�2��*��&�)�]Zf�Yec���Z��)�)��Q*��l��v�C���m12@ƛ��*,¥Ah�<S��g[hu����L��'>B/��N�BG���U�û�U(�Og������k�-�ѯ�!s]�y9��Ay#��;[���D�%�ݹ�I*,r���He��@����^F	4kR��UGNQ�˛�;_I5����Ƃ<ߺ�-�VO|dt��m�ak�-��:v�	$�vP"� �sxx�'�����������cF&��6Jy�Z��He��)"�[+![�u��-���Zh�:zt�B���{%�3�FZ�h�Ң�EX�
.æ��<�	!�t�5bKg\�se�!?U�ɴ'�x�� X� �)�Q��(�M�KP�i�Q��6�R���P;Y�h;�T��x�P��!�D��V��R����`
�<n����CM&H�7�������A�«=��G������ �xk��,R��@G��x��;⣁p�D�x/�+D*"����o1�z�y��=m��u��E���2��+6�KK�A�}����!\����_���] K��K��7I�r	]-}4�B���č��0"���|��������w|��T-��]Dg0�I�ޥ"Wf�1U���Y���4�Uo.�nX�ͯ|f1<{�8*�ln}�?o|�1O}V�Oo�׸���8����+	*�]Y�����H�q"���.�|7�P7��Ӹ�H$x�y��wF�ѱ���7����J���TMt�zX,YAz�qx��ӓ�K�p|���;�`�ot��k}���>�Χ��5�K�����H6'm�� \!�Ѳ�l`C��^[�j��ۏ;�m/��;Uj��Q�q�{��«��/��N����x�T7#1��=�G��n�I"_0+����S3��\�t�an�j6{Z��a�k�c��l�\��G,�mm���cWk`�~t�l����\_���#&�m�{��ՉQ�0���|��{�����9b�]�[|li���MϞ �:�nlR�bQ�2�N�q��t�����O�������Iy��+�F�ע�4*6�M,��ױ6���'M>>�[A���_�l������n��7i�=�9��c��UU�i����-}><���WG�ե1g�۠�[�p�f�����_߽�}".A=���
�[��1�����L׳_S��� L�S���a<|���s�I�=��k�[��D��<Olk{4�6��������,eŀf�Ҷ��ms�&|��6Mnuf�-�a���©�kٍ�O�����MN��/���\��'��*�������{�x����2!N&���
T�:���N�ډ�
��X�'��P��H�JJ��f��<��ϛ�U�CJD��,1���UM=g�p�Y����Rs�yga�X�dTM��m�ʙU<�8�%�FR�<qܓ���xilB�!� �?� 9�Xb�pbgSJ��ari�EϑG]/��,M%rjd�"&#�i�Ә�Im�>��T�[�N-$����}�l�i~�����5,��V���Y��k�u�$sA!���ZR�m�57����:D* ��|r�V�?YsS/�P��]������\���E�R��SW��4�|$�pN!��Ał��k
2���1���-��P�'�9�����F\�̱��`�rȝE����j5,E���^�U�2� 9��@����7��PD�D�o�˱����g����ko�s�zZ<�f��F�R�:q:Z~1U��,3���@�u ^��`)㊪��L�NMh��R��Ɋ��m9%�.Pu�j��*+�7�o��k�h�dmWK8'.�8�����������|~|t�}+��5˦�W��f�F�������k[�O�g[\�1�_�l\-�k��-�`;��r�rƽl�m��MmlPDt��J�`�F��7^�j�ܦ�_�v�4a�$�[�s��-����`�_>��$����Xč��o�<	�ƣ�/��w����G�������[i��#n�o�'x��?m�s-�;� �[}߆�s����'.n�Ir�o��:u�,<p�xo�eЛ[�����E��il|��7��ݕ�[UVV�R�هI+cc��x�X��?-OB\j�%�e�A�4�=�y�f��*Xyۿ��b��aK���������.����{_�l��67��°���B���7[]G����Ac�ߙ  r��t��
56�-G;��QsH^�e���RIa�����,Q)�i8�(ϗ�30>=?#�'xڠS���K�A"�HU����	�{~��1�� ���a����S�V����槬}��Es�Ԓ�,zXI���+S���i U6!ղ����孛0�y!I��N\�?f�cr0�c`��	ّc�f��3�7�[Q�4�u�Dӱ�[�(�cR�J��`�dG9A9c�3�����&SS&3r
�������h!)� �� ,n~^>?F*���Ş%R���*�ǐ�a㌔ՍV�+�3SI�џ�`��[L����|z�o˥w2L��ӹ� �q��Z;���ac)9�k"�/���]�7��!WC����i�d�$F��	 t'k�$�zEŒH�A�����)VN̬��4al
�'RՕH���|���mmK�&��،iu�S����[�]WU�k�#c��_��S9{��܄͛�7ۇ��ʧ(�e}� �/���æ�_�lk{`�.|ͷ����if���ƃl�<k����k|��~�������.J���lb?:As�V��gM�����B;�w��\~|��g����s�q�m{������Ƙ׸6񿇖uՕ��
>_i�x�����_�ֺ����_�� {�4�sG�l4���I�\X��pz�m�a��� ;�5�-����������������k�������7n��p#�m����x�uo��,����I�O�/��fv����x��.	�-�~���Ƹ?q� �K�l�;��r����Kj/�j�Q3@�sZD��뙤U�t�|��ѭ��-����7�C�]4�^���M0n�9���	z���̮~�u1%�v:����� p�r�L�Y��ݣy����I��%��(>�����mN?'�~k�J�XVx��*��9{�J�;b��R�^��Ơ}��vo�!mM��,��3y�e�\�3��0�EvB��v̺�lm����Nh
�� �����ݏGꢩ��� n���� � ��$h��4Z\�k�X�C����_��/J�`�<���^I�V�<����$�kʹ:s_�av������ ��1����8�1"��|�$_�s�QQ�tԎB#Q����%�7��|E��8V�MF��u�1a��h�/b���[vŀ�>$m�}�o�� "<1���],�a�7���[�����ܸ�*.n�F�g���)R7=��~��}��2�o�#2{��e��P|w���Ys{M~�rS���lI����f�[�����L]v#}6��)�c������ ?����W.l絯��O��l��c-�'�o�]���.qsa?Θ��[ko+����o����%D͕�(XGpr�P�J��}E�醈�ea�t����{]��E�s���襲�os���1c�ÿ�=����Nt9|��>D_���_b���>�2�`�c؁�ǽ���t���*5R�2A�0���e(zXt2�m
�m噸�tPJYR:yd�.A�"���7�b1Q-L�G�����]��w��Mm5`F��;��()]���SSKQbޮ����-t[���}�]�覩^'CF�Ag�|� �2�D2�UF���l��Ko��:� �� �hq���� �/��R-�IIN�~�hP��^؀@%QE�#�d�B�gOT9�bT�&�ROH���9q�v��_���d���a�)�ݷ����g27��t�om��8�i�b*�-Dk�R'�y"�,�u�.�eC���Yě�����E-�;j�$�6wc���f�DLJ����~u������/���ig��GW���^�F1�?.E����s6*�
#�I�h�yC|���m�0��*�"EX���{��k}#�D��\*�._P<��E�����cs�� ��0�$H�.�e��sc���\[m6Ɨ6����^��LxxL6��xa�Q#��[�����li�#m�� �>G�=�DK�r�.��غ������c޹��n�77v��o�����Ӿ$`57���|����z���-��#��YS<d�Q"ot��2���R;뿖ee6ͽ��n9�����#����~X+�R<mo��f	�l��_�|5������"�8��]� �/�:���VП<H� ,y]��M�k|H���5H9[+G~�u�kwB7mm��2*����m��8s"9J�3V��9m�.�m�� �����6��:b���ә�/�JZ�A��z��B������̚�3,�Nul�hфjOH9۪�ٜr�}6�z_:�H�/TAp�@����e��u;[���d�fa�c�<�"3x}⚲��:ک9�**DcF岢���nY�`�̇\��k�#-/����p�*������rfwʺ*��9����x}���w���tECWP/����ۄfr(��Pe���B�B^��u8H�"6��E�k��H�,4��[8�+쪠�[S����]� ��.�C�`>n#�hd�,��ݾ�F�������>ed�X�r�fN��5��{`*�$2����{���m�mm��>x���Ԓڪ���l��zx�� �=� ����\ph�H���W���9��&���6:$>�
(��tL�N�1,���J�@�ˑ?��L�IY\\��a���ap7�q��B3z�Au����ok�Lf�����o�[

��,_���'���<� � /����êkʌ� ^�[O#�ƺ��`_Q��� ��س�F�?��|qo��/��w�6팶�}�A�1�� �|�k �������M��цko#�嵷�4r�oUNZ�B�˥��Gm���{^2�sq����j�_���X��>F�����'7�$���'��]]��o�M�MDi�:hش��KX� ��l:��F�|p$�al�]Jخ`�.6Ͽ��~N7����	-�o��a����� _$��pW�؝��qs���A�9�W8+������;���co������f��5Վ���t��>a�?}����<qc��p�=-�f7��η���Q�6h�h�t�� �;f��q��V~�Zl������<q�ٳkC:�ϭ�r����ڏp����iܛ�5��Lgc�����y_s��т�1R�m�ψ��~�e�ݖ�G��{h?;~�5R�,t�����M�9L'�p٠��G�]�����i���]A�:�Am�w��_tk��Ff�VC��3��.��՚�x���)���!S�wfk�{���t��2�\�����a�8��gf
U���hA�0�IL�-nh�H���mҢ�6���r��TQeD �����B�d�6_<�֪��?�=Q��ऩ���&�~�d���g�W�Uk������M����C�8��L�����C�X��>����k����	�����>�#cn�uH�o���卷 ���	� L1c��l�#�� ?���w7��~�X_&F�ǔ3������6߷�����||�Yؑ���� �v�|]H�Q},t�Ͽ�.�_���1o?��b�;�^�^���|���:y3�/�
���bõ�d]u ��\~�7�K	�������1o���6�lh�w8�l�[���V��>8���q��*��U,���@��!�a��`í�uX\��()�t)(!ݒbR��'ni��/!)*!��"!H	�Q2`��f1>���u�s����羏!2b�w�g#:Q@����I���29 �r�w�I��t���P��)���#�T��l�R�eT�s�/�Yi�9
MLὨ�1��P�"w=^d�C>[����-�ɥqkV������ݏ^U��ه������)��c��/�=���q�tQF��L�B���������;wz!QF�[a^"e�7�/{�4��a�Y�v�� ��Eb�Y��י��֛���f4��?%-��}��)��OzS�0?�k*�w�
3��ѷ���tXW��C�]���n��!�o��f���O�������*l۾�[V�T���M�%�S�r�f��QU^�H��g�^`Ҍ�^F�]�����UI�~'�}2&QSPWP���[鑚�﨟�Lw����Mf�6�(G<I�k� L��'�xV=L�Q�K���{�f�[�18i�+S�MSF�Dp�9��!k)�48)I��a.�0�܄�DZ�B�.�<�4L$���&��w�k�dh,�7�?,c���O���:@?z�Z��M_ 
b����t|�ǩ�a,���� ��쥴�E4i�|�B�Q��ѧ��p��S��N�]rA+'��7��A�h�v���鴾	�/�;�'"�[��O`�3��MO��̄�����i�}�N9Oо�����=����:�U  ����/��E���@������*h!� ���},2��dOv+��1��d_i�ɷ����� )z ��K���o�4E��ʫ����~[���n[~|��g�{�/[
��ŵHVp��ף`����M�<�?��2oh������?@+�����m9Mŕ�=�q��z��4�E�^�k���v &5��D%���Q�[׾�oM,�"8-t�7��,�}Y���{26=+f�t�&��[K.¥�2��w�Dt��,ZBWkk>?��,��j�8\||[Yq�o)�|6�}�ӛ:��Q�M�M[�}xB?��R�c�j��ɻ"����I�5���ɮ����ʈO?���O2O�5ʰ��m-5W[��61f���]3_�wyG�<�F�ס�N<[�Y��i%n�-�,���]����� �{Q�KFݸ�}mS�앯�G	�9�Л~����h~���:TK���C>m;��L��f���k���D����O�����	����~
`�o��g�~�t9�Drj������0<�ɐ�)�V�Z��FѶ� \K��55�1��t������˜�Ě/��Ю��1�OX#@|�������D� lsofMD#S��5�uN�'��cVi?X���W�����n��>KP��t7��Υu�u�����Nw�����w&�wu��Δ;�[�Z�AB��2 {��yD=VzJ�҅Ǵ���[���\E�h"�|�M��S�����W)�Pr�T׬��(�����\��N)7ƈ7Y�&7q��z5�7�y`�ggu0V�p�����]���Hxz����Ф�a��tbm�LNږsg������!c2;R�B�X#�CB'b�0#Ķ���!�����{��0�'�J�a]��0ꍊ�?�X%�:����҃+?�����&��T���f5���G��H�*�Gm��\�t) b��l+���;{]ixzr��l�K���=�ܫ�������T'��.�M����۾�/ �!�H�g��L���m<
��v���O��K����N���N�h|�T�w'�-�?xb��N4��-f��8�,��x����:֨4��wh0	L��.�|-s��G)>{��)���V���D��B����_D9]��5�=�x>]���nbtY�����[�������'ksGgl�:������_Rx#��>:��Rt��T<zY�t���
��X�z'�zl�5�5� �$u�8�ާ5U���x_:��J��,zUUy�p��q����Y]��Gő�;E_m,�'���Fվ�%$���?���A,<�>�������{�CSՍ{(���hI-��[7�Ђ�mcz��~?�q.	&Vs�u'�M���k���u�`�%+������w��^��z��x��<����dF
-ӑ-��Ɲ���fd��|�i��#
:��{(��v���ocA��M&�1�!�֝��Ƞ��^ᦌ!"�2����]�����7�\�G�R��B]�L�JQ�l#�3~�H�i�6�zU���%��+���s�&�`}�-�'��NY	��rm1@J?RSi�࠳V"�MR�~�]<KFp���U���0Ox:&�ϒ���ě��q�x��N��"�x�J9�[�;�
	�F"��ݦ&}K����)T�&ht����s�F
�4����	�J�cjH�)�Jz��"�C~4I���Y�~uh���}@��	���/C�8r��m,�e�'z����� ���(O�v��k���'ݤL�`͛�x�(�y�&5���rҿ�Ev�D{�:��G�`!�Ta�r��5M��Agu���. �X�18��՛<	aڤϳEN�}TK�[e�Y:��UL2Gk�����a,|2�&����t��&��wtAA�Ɵ�z�#�2طj��]�^���)�u�z�9{Z
��'[�\��v�4���'z����ߣ(��I�u�o��&����ˠ���ԃK����hj�*�Q�)���ܓK33��<��(�Ƒ�C��Zj'���n����S�'G�H/`��lM�TU��[�E���jfPL� ��s��uq�vǒSfp� ��`�d����7!N�߲��?YJ��p[�$5�M�I��y�oY��ջ�����2x����~�f�y9Ņ�,�Ǝ'�a���nw�D�&D{J��)j�w�VPoS�m��k�&�]&�%�-v��Č����ԣ,0����(~/b����s�u�%��]�MQ���U����l&v�c�#��[��R5���4>��@������ثz ��u��ƆY �I/�S���&���W�ԇD9�f8�I�1؝����3P��|�A�B5.0�H(q�����s՝�Z�~�١�̞��H��� ���v�-p$��5F폠E�LՌcj�qOj�ي�?���V���2�	���ԕS�E.Ó�@>��+X�ݝ�X�i&�#D�����dc�����G��+r9�s|�,�)$E7|���z�����g����Q�x��~jo���Q�y�c����t�N�tu���>"��֏(��1��^��S��vK�YU��۪�]��� �g���m�S���������d��� m���W�)� �:�����S�ڌ��~�-F��P@�T��C[���;��Uq4B
��C|,�]�f�iM����?�?k��լ%&&�a�/�ù��"��'n���n`����y����z+����3���9�&��|�g�w�&�W_e\q;�nԶ//p���Q�5M�|�ƀ�ZMTa�_�V۝���\��r<�;����^}����-:M�O.�/:x�Mh
%��4�&��L��^�����H�׫�Ð��ؓV<#?i��I���dBG� aG�E�wm)�T��i7{\׼̝
o���e �����ӑ��������e��I#q%K�.�n�q��M�������wV.~zi����}ġ��`����}_<���B��&n\Wa��������v���A��1�&��6+&H�����q�����]9��b7�#d;�����mn���8����2��N�a�A�7C��	��2;/7@#k�'��t7M>���(&�q���]/����׽
Uf��5?v#���j���;�X�A��W�~=vԦa �����1]�뎵��۬
QP.sH;�)��˭�~�K��Q����y-��1n���% �uu�=�i������>$�  ���tt�i�f@���O��YYO���v2�I��^1n�m�p�Tyo,ZG�Y�݃]���=���\ t�v"/ �;/)���&�\ >�8L�w�.	��;�v� H�@�K��p������-����t�}�?7\s\��f)te���|
�պ|�a��f�aIU&�/�9��D��ۀ_b؄�W�>~��+$zQ�f�>�o&���F%�ݡ��7Z٪�]���E[P(,{��x����$��]1���|���Ѕ�h!\�z�Y؊�Xckh|�+H ��J��_4T��������ճ=���+�%�X�Ư��"���~����7�W���������kG����̡]1�y:-������0��Ek��{�%kV[� f��<-�FGģY��d��V������޹�.�7@r��`�����ʐ߸ȶ�6҆Y	��fh�B$-%Go�KΩ[L�S
h�^�� bz"=T�4����7��������;j�. s����n��Q��ŧ�:��S2H̡�u�`��owجI���a#�=\M}A�Q���)�nk�=���er�É��R���B�6���}1�%��߭�)�-ʤ���ɰöԙ׺3 c�šǘN������� ��-���82�j��Bck�@ؙ<�_H̕�/ۈGV�C�%�"�g���X�C��3M��
��©x$g:¹y�חqr����ODl�'ۓ�d�t���9i�������=5ڭ�?�EG5.'C�~�����R���s���9)7Ef���5��GM���ĝ���~�:�?��4=B��O�dS�Fp�?��_�R��M؆0�}LK��k�Y�W3��9�:R^e��$���21J�F��s~��`�6ù��>�*�����WI�|9<��w��N"�=��D:�7�B�@���o�`�g�8��Y���w���/���,��A��:�7s>ʺ'xɴUٸ��.Nݦ@d���D����4���O8	W�G��`��6n�ǥ�� ��T�O���	����Qf�qn]�OoA����&^۹��R}����OSe���������(����~�Q[��y�"o��d5�Q����N!>m��^�ԫj(�48��Ka�%0��r�9|����̪t��p��a�*�s 8��|
���Co�^���Dܢ���b�e���?�H���2b��WDv��$h� ��u��P\Z{�ҥ�g�P�����~O�Y�P\�� B���2C��ʇ�E�勩S��#čo�3L�W�6�#�\L�r`�M��X^���2���:ʛ��E3{��U�ۏ�����������{�,7��?��7�P�6H5��,�����.�B7�tl)��2s�u�-Xr-M�z�ib��F���L�[��A3i��/��:�YU�;�5�'���0Q���<I\||g:��aR~�m�ig���1���w�s�/  ��r�:]�Y�.$�/-9���m�Cry�=Gȫ+o�9y�lp�2����<��|d;3ݘ�_(qJ�9>gZ�e�~�DTv�@�����T}ճ���zm|�a���_���z�28x�((,s���G���Z{��i��z'5��E@A)��u��zLʿ&�q���~���
�������Nz�D�`�w���Jd�CͽW��D��$ߨH8]ϸ��G��\I̪���*W;�L�*+?EWM:"�-|H��:���M�_�����\MT
w7:�P���̏vf��o3*"�F����Ogf
�8^ߞ-�)�㒲����1L`�T���neW��H�K��Pt��3�Z��w,c����8�O>6�Ͼɉ�"�@�X޼��PX}&�l: 3�x�����Uޟ� ���%S<��z��rbZ��r�F�B�x5z���"��Qw���1�A�����ж��h� �������. H�I��-<o�����A�	:#�>=S��Z�N��l�ۖ%���k{mç����;���d6��<|F��aXAD��w"�h��;ɪ���:C,i�Y��$X��K�<��g�Sg�@�JH��{��Se�5��n$w_�SU����wW�a�cת�`ңn*O�V�C��18�,����}9qU���ߋr��׊|�J�j,<L����}�J������#ՁN�:���fF��}�_NR�!m����|�r��ͮ!��R9=��s�4I�ԙ��ۭb/���*,�M�{ǳ��G������w�F�a��CwM<�؞IFiM��	�������X�\��`r���A����x�P�y�������u��)ʏ�uP|�U]��o>5� bv���A�X?����>��1%���T9�1z�ϓĹ��Z��7@��G�P�g�fs|u:�80�f���v�kwk~iM�ֹ�<���?�����х�翧t�l���&�_��KC�t:�R̯1����ok��u���M�W_L5�u�������}�)4����qF?ޢ�zi��(C��g��~��ΑR��0��ΉS���Q�<�ik��(x��NWL99,���[����ݛ�v`p��|.T��/&Da3UG���+�����YKjSΒh���jSa�s�BR��?t�.�nE.�:��"J��6mK�|ʩM��~-2��V���\� Cb��2��5.2��ݷj$..�����&~x�^ω۩l,ݱ:�D�w*�5t�����d���5
Y�IF���2��5f�)����Q<�c�eri�WFb█~��?�����@�3��E�J�,�<4NO���8�����r<��`��1-��V����.��5C;�Π�m�'1�o92�ՇH��~���w�IdE�� ���j{�&����r)(���C��*��#��+���ir���IUnuK�'�=23�#4,6o(f�9A
�'\��W�bl{�>d8:9z,���V����uv�x̠�D�~��֯��e�5<�v7�nH,�j�k��.��ކۏ��.�N5���䪶���VxOҥI�w�;)��N���U�E�>�yU���E���4�7^��'�z:V�E��(O^:���8!�AA��K�ϰ	؍�e���<���Hx^U�_�*(A�f���L���8�"�F
��R��n|JUj1ȳ������������w��� 7��4�G��:=�x��?�l��ӚTD[rB��]��PY$�qE�����tI�!��lZe��J�yt���pu�$�Uv�[I��>�WN��Օ�_�*�y@�	KF�3d��4�ҷ�]�K8~!�J�g!�0��U)�_�Zl[B��:�Yӓ�<�iB�N}�m�L�|�~�󳮾m����m6����	 ���F� Q�Zg�)
��>`��T,��.���&F�.�'.����z�����7�!����Bi@`�K�sBB��x�M��HA�/��v�������
�+`frb���4�͞P�$� h#�������l�h����T2&�ǻg;���_\�z�����צ���| ��&"%�Wl?�Hy�b�ش,���:����W(S��SX��+c4�ag���Vڃc"��gO+��]_8P���(���ڻF�ݑ*x����Nq�C׹���H=͝��O���?���E�#�+�d$����a85x�cy �ES���c}s�B|";������+ �ոS��l�KJ���}Y\�[�P2��]�bsm�2`*�����o�ӵ�E��z���z&�Kы��ʦ�k�ع�6�?�e5�:��$�d�v��cc����&�`->�R���㵉�EAQ\l�ѯ�~I#��ʩ?n��o��-7���c!���8�s�0{���X���n�"qnW����'P����|�7���6~�D�O򟉭� �5K��S����Op��ݔ9{e*�h���S��UC�7x�ص���KI�w\j\��MU����nT���w[܅�ވ��j�JE��b���ɞ=��;���� �u����$o풷�00C�x�A�$�8;tz�I�b��T~��A� ��~�ߏ����� �\p��׾C�k����<��T)�`.�V�ckP����g�*Hp �y������9���32?9*ԋg�ٝ�b��3%��-$K'�$+��1�S},"�z}�!檘��a�aU��12C[��C���qXx�ݏ�#:��=TF	8��}��|�֢P�8ۄJ�ß�F���yR>�x�u���w�m�M����`k3<�w���{sR�kD �S9��W���%n�Yb����[	�+��7k�����s� <�<QB�5����T�p!ųy�Z�g��!�)����T[��~I�x%�]�T"�[%M���z:���w�	t<,�߶���C�[�����V�܇%�|�~+��Iq@=�j'P�����x�-�8�fE[�Ǌ#���٧K}���n�p�}��Q���{���L�a��_��~��D���N�:1 V�b\������џ�߆�~k����̓?���~�=�u.�drnh�M(TXE����PQ�𛯰�����Q��+�U�V��bjv%��O�#LX;�9}���u���~��WN<�1㡛�?Y���
V�x!S�AB��|+��˪�[w�I�/�TT�ߵ�XY^j��d���}6�+�ds҇+�P����Ocm�=	���wM�y����pd��X��Rly5������W�l���#w5^���d}D(�{z����	.3�:%{�h�YY�F�[�ݺ;�`�@B6�@�g�w{

�OA�(�-L��wֆJ��EJE��V��^���Q��:�y[�tR=*E��"��t�<�!.�=��������tt���� �R,1�[a���9s>�(~��lr��I�k
9����d����^��l��s�*�O1�Qm�H�K�V��B�rA����w5cs���p���-�������(o�Ƹ�u�n���e����((��)�A@�ߧ�����Jt&�`4�Lᵤ`$�~U�c�_��<z�N�H�=�W_炚�9g��n5j�o�+��!�#�#������)��Id6�j�1�;��1��b�PuL�/P��^MN���P�a�+���c������B�����d�|� �,���$w�
����x�������%��Sj�f�ZG
ВR����*�oT�TV�V�W>>}����Q��]C�F�*�~�jèS}Đ�Ve7��a:���q��2o����0ۿ�9�]�K�JN����:�kԻ��H�Q
��ѧ�V�"���R?F����D����?�[u�,57�/���d�x��D�끳½�}u��)wn0$W�˶��ǔ�Ǽ�{O��/�0��d���܇*Ko×�$��,�§���o5մ�4���`�}W�s�b֓G߆�|�_N}yw�Β1h��5!�M��0��Ii;q��رƂ��%�L��s�p5�9yS!�r�!���&e}����y6���p����D&�S�=%�O�z��T`-r�V|���O�R�p�m��!`e�P�O�A�w��0�<8��g�����Q\]�?�Ւ���4c\�g�`>�=^�@�L(\m��9��yy��(h�Й�(p��|6�f<��qm��G�ٔ�+a�PƩb�<���?f�n�X0���O�/��Qa��0�����^G���`�p���Ap؃�'���tSS&��R~�{w'�D:;}��hr��g��dy������%y�𔶭:Zl$'��)��?��ѯ�w�_s64^ ��a1�'����/����*���_�jk�)<,�JVq1]#E�EV^�ZG֏3}���_���v�#�bf�%�>���!����K�56m�u�b��O�$�zlN����'�t�9j. �	�dō"��8���R">D�^�봑tH�%�?�Ҙ���,�f7�@nX�@�9�xt�����?���>-������>)Hky�f���/�d�n���o�!8Z��ʞ%5)����x`0�c�J!Q6	FѾL��ս]�-ѷ�+i��XP*-�uy���`�,ƨ5����qd߿�OS���Ê%U)+"�Ư��U�����V��}���3�Ű���(^V<�ܡ�5G���w�][ ���8�&��3St�?8�Q`�����S�g{-� 4t@Z<� <��lҠ�g��A��LM[��3/��q���L�h�7������!�n�Z}[����>�	���\�Vg����:���j]ˑ��\�B�ʻ]|e̓��{H�Y;[z��e�M� �"r8'H� �|Ј�$cj3�b�:��;���C�(�i$k�!/H��4�	>����W4,����Ĉ����~�aϏ�!��H�D/b,�{�ާ����3}�=�Ӂ1A3B��M�t��J�⩉����=�f�|�4-��M���&jce��b�E#��@��Ͻ�u�e�7���0e��ܜ�	-��dߩ���s���q�	��7=�x�V�8���GrL �{��
�[]7u��
��-q��p�=ň/ �Pt�sT�ES�:��v^�`S���'.�������U�W�Q|����9F�'�e��_�S�oF�~Is��X}3�����z�;���xF��@����)�*�`e(��u�����&�k 5T��#�Sʳr��C��?@�=�畿�*[3$��x��r�pS&4����٬�;KL�߇?ʉ9�}&/�-\�a�W������]�F$�c�:^����t>�5if<��i��}����fy&-�ޤƟ���o>�z��-ӥȯQ����)���T
x]|���v���&��H��[���g��{x�q��T)gq��s���֣λ�����v'�[�'9<��\��O��A���Fp������E�ݿ��k*�y�$��F������u���"T !��+<��ߙ(|44'� �K�W����%�Hk��pX]
��N?���?��q���z;iR���M&u����Y~�{,"��r4:MNx����U=� �R5\v<D©!n��P��B�aÈw~�7_��]?���ˁԟB��F;q�n�}������ϻg��d�����S�{*XQ����N�{!�j�^�I�_m*l������<e�:��Bk[��IB^:����^"?���v�߹ ��?���b�W�zw.��&<�egy����}���j�/`Vý>w8�/'9h͚=v��>�hǚ6��8��{��[�D{�Ի��$?�wM0��1�Y��;	u+�+��xϥލ]�V��3fbQ�
Yp{�R.nEԮ&��XX�du�g	�w^��e�(T�V���^|�q�Z��P�s@��2�['Z��.7��*��i��7�-��߉W�<)�	;�`orydxKw۸�*UQ��'�}��g�� ��\����PY��4��L�G���9m�rr�"fֱ���������������+��x�U�u��]��S~ŀ|[�'�T��(x���J�6��� 0s\�}!��
v3\�oPdv.�c
��v"L�E:�w^�)��)c�qpWN�`�OT��&��µ~�qNSS���L�څ�Q���9�ʵ�1r�f{�I��(jm�"�D���H�N���v%��Y �@{��d�r��ۚd�<����i�_��)��[�~x�`O�ar�|iqED,|��L}~-��^�(�����a�& R���*1o���0����1����z�"��ޗ�-X��;�Y�u�eK���Q4b�����W�Y�]����,K�y�
��� C����S�# ������)�3f�H,�|�O�l@5��9��KWml�9:��\�|D[���.0���h�[?�R� ���z��wTi��@Rߜt���>
	�����~��V���VB����z�1��>w���NG�3Ԟm�w@��
ۉ���ˁa�f�[��Z�G� �	�vS�	���w��3	�q@�J�w�1�tt��3VKrc{5���[��Di�~���v��6ƪ%9���%9 WQ� �7c����!�����Չ���E�)��P�#JS�I�z^����cӹP���_�Ъg����=c�g{E�D�R��Ǝ�2�j��Ԑ1Pa'(1�P��r|��!țt/\�PM�O��I0�W����Q>�-cCH����?��C\��'!��h
uJ����0�G1�X��~4r/���0�+���d��Ǧq;�ؐ��K	'����{�t�R�(�����>a��<��@O&����>��ء����H�V��H,t��g3��l��Z��C�x�p���Vp��1�����v]?3��B��#��� N�2�s.�Ip�+����q����q	�!���w9� ��)�Y}�y�L쉖3>�>�A��)׿]c�x5�	\y�%����Eh��f�Y_�wzA��a�x�-�#�Ĩ���[^����&�ؑ<�a��'��"k^O��oe&�ۂy2sݤ��n'�'�/������"e�K]o|�:��=�$͛��-�w7ͅ镬����~�	�;�?��~��f�U�����N����UA�����ж��	"�7�����F��Alz$����	����a��F�ͽP�3d�������?�Ξ='�D����|����7� Tg'�͖��=�����C�O&>ryQ�9E� �i��b�rh
*"�h:�;}Z sR��&��1��!�{=h���}!6��f+�AOA�)l��jd��Qv��B����!�q�{J����Rt|y��0�)��kTa)�Pk��4`�K�
j�#���v�q���T��>�τ��\DCc5�B�����ڣ�)m%�⃺"��ᄍ����6������s���c���x�f��f��C��67�ݔ�Β!�[<x����б`���L	� 4�r��� �d�cj�1�,��.�O�O�N0�;��l�c�s'-U��F�I����K��������=}3I�BC^��
3YG��*��z�̯��u� �����>��ޙ���EG���d���:6s��KI�+���:+w]Y���(5��O�۩�	A�b=�uQAv:X�>b������v���-�ĬR�|��Ҕ��M]2���3��+( �������Q�܇�c�����땫a����%���Y�l���LP?��u��i����NX�12��R�w�|]�TI��٤���O-~��\-5<R��mڜP��e�����D�������=1�]�zc]��i^m"[у��#pV��!~����� �(M�>N���h�i�V�TH=�`Q��'�5m�eE8�L��m�DR)t�	�n;�7��Ա�Z��W�Ƕ���qy��LXN�Om-'saBA�:�� 
eq�V@?�X���{w-^��)*�'���6��������K7����tu� ��	�1�A�'�!j6R�Q�-Dհ$�V��ֹ\��q�.� Cv,����9Gj�K�\ f�1qH��fJ k���@^�b��<&�n�mT�x2-����ص4�~�ɥN3S��1{�Wo�:�`D�a֜���R�gKP�~Yw>o%�Գ��@?��f[.92�����(�����ѫ7���G����|�>	em�Я-�����?�̽2}�����O�r�t��x���NCc,d��[�m�`}�ubV�6ޝA�y�"�msק9��h����4*Ct4h�*pW,���1���XS�C���G.��a�SFf�-�&�%�nTe��43�-����sS�0�|i��ҝ)ݽkt�������q��@<a]"�Pv���f�J��_$8�
X3���q���X�Ěu�(}���)���4c����\��H�'�϶`5:��l�>�z�"������I�)�� &�����*��!������x���)�-��Z]�\��Fຟ}�&�I�O��:w6���v�n���
iz�:Q���o�����ҶY��؃k�5�m��K��I�y�R�N:���
*�0�4b� �׻*$lw�x�B��V�� 笕�0-���3��B�W�fH�cj�������M]�WJ�����cb=|d�/�>uH��Eq����$os�d���骨�O/p�T��3���R���%�E�w0z�m�(��z�잫�M`��8�����OVl9���ΧO�^+B'�"�y�M��=dG��.�w����^a��[lFE��ˁ��n�އ���}Z�V��L�xS2RL��Wd�����W����7�1��5���;����%+r��x�^`L�d�K����ҧ��S��OZ��<�p���L-��q���Pa���-7,��n� �캐��X��yE��Ǫ�J��k�Q517�d?u�F�+?g�)K��7��~��>$���[C�k������f=��x��������x �@dy�y����Oӆx����*�n^EQp0��C��	�����k��%$�^���� Ex���+ݩ�(��k��C���h\y�����x�O��D~I��#>H���k��-ol�̸�{�����-
^�Y.	�	,,����!���Q�=���Z�.�?N��7�	�ȯ�O���q�Pv����y������wԟ�N�� T�ae#���5��sqZ�qHh�0t�o<%;Yz5�8�s���������o��88��Z�(��%����r�ڛ
։�WW��No�w���ٮi����W�|L�5b��X.��&C�L��;'�+ʐ��|F�ɵ�����D��B���LmM�b������kX�￨�ɓ�1&�7��>E���.��,uMK�ף��+��hM�J-å��٘�Fe-�0�ݥQ��R�|S���0S Ro�6lz��k���'ώt������ֿ����I��Ҽ���=�f)FWr>�;��q�PJ�1�4�[��-`�q�h���g(
�9�͵�(?-����l����r�I�"�����U]r�i�U|�"9���\I��_ɦ[���m��S9L����Vྎ���\���݄|}&܈�Rc|����)��rU���%@AeC�5)�n/ї%��Rw3�]��#����S�s�x�5d*�*z���YU׭�Y2IBE�ިNI��胴���n�-������'��k}B�Ʃك�����a]���a�&�L��P�b����w���9��cg�hP����������IW�(�.eoLb\���%d��q�L��q�t]�P�6����rz�|�#;�a�Dk��N��嗚����;�%^�/�?j�X��4,�ab��΢����w0�]Ray����׶F��$��-pG���#���\��̓�X��K����s�B�7�Oe�û�q�y�L��o�ɯqhI�v=ʘ���O�j%ⴴPt��0�o�g@�6�Vm�	���3���f�������������SX
��I#�?�ٍQ�Fg��j��6;�ipq��
@��ҝ�Gfb�=����9!! FP��F|�w�d����RR�&�|�Ӊ��.��-n�k�A��-��f�xZws���#��批mn��6��0~�Cй`5�m��-&����%n�\ �b����c~�.j�R�RONS�� �T	X�s>�e���EY����g�B8So�)�r�~.���#���>WN���n�!����@L9Ҏ�Xj·92�N��`VV��7O��oTUn�&3"Q'��{j!�($вv��4�_�GU�fO[/ YCw�����Ίo֣���V�z
�r{D��|�Z�X�{l���1Rf�|"H$�7;m�~Ny��g��������\���r��]�tk� �`�R˜%�9�/jIRSU~�A��L�e@w�	+"L~l���TMW�g�����?^��h�h�-p�����*9f�R@7��ug��;~+��A�j润��z*�jq�,wJ2|��I�G��̀�M{�����-�2�p_��R�L��pK͌�v�B�N���G�tVk~��]9�B�l,�0��T������/�WF����*ܭ�콊�_^C�&�$���41�
���c���I������:A$� ��k}e���#���R� ����w���ApŬ�H��� �U��sY~m`��p���+�d0,���Z}(�mN!|�bLD�}�� ��OU�f|�:4���nd������觝!Z��[c���F40�R�������"y���;JR�B��mZ��̯ܗ:vowʷ'-�5Y����Uc!6~�!��&a��M)}7���T�<.��JG�	w��`����0X[��_���	o4/�	%!O曁t{�����[<�p��5Xׇh;�w��J��R��<z�tX|��pq8r 4!��*�W�Tȃ�T�&R˙��%��R�l��3\�O�p�������B�>o�B���/�p��[br�F�
�����{�EA���%��T��`�+κ��6V��C�� ���������n�_ˋ^��j�%�XN����&�K�w���0�^$NU�탱�����g��'�ڂ h���'�����@-�pF*��WzO�? N@��s	ch�dWV�Y\�V�n**�|�d�)#Nc�o�6���J.�}�nra�����"�a&k���7|�A�I�f��:�u.�R�N�mc�:��|�H�+RL[9J��hf�r� �������q�"h_4|>��Қ5?G�&1��:�^��ya�����}����� Li���^�v�ys�)�jܻ[):�U�~�ْ, �P�`�r��0���w���H��,A��?�5 ��� </P������X��$��xh~�d9r{�PF�������v�v�Mwa� ��6�>`���K}��Ŏ�= ����/q��F������S�~� 玑���R4��=�.�Y�l?������A�Z���Ğ�����yF�ť��L<�\v����o���6��|�~�;}�^���y���ӷ��mp]K�����`�����f.�c}[ůn|D[��C[_��������)��.`t�D�ŮH�:��[V�̧kjT�#n��C��CP�?�m 6���M��a��]�Ռ������k���Tٜfes�@-g ��w���m8�KM�^8�{n\��왈�cˏ8�V1�Z��;ފ��I�OێO08_�X���E���.Kyc�A��ն���g]�����dS�o�#������o���+�"�*<��������\Z��1]M*�TD��N "���'����<����\�p�wR��(�bƖ"K\����&6|�Y�kj��M6�e;�����p���?�)����eHc2]S3�cm�lN�Zɽ���&Y��
�D�����5��Y~� I&<��a���$R�9$�E7�ȍpYh3(6�*(�kw��>�n��[�r��J�5l�J�[�6c��7�r�ݔZ�$�2��N�-�$KYcm�� 7b��_7O����{�`u�k����7���V����������� ��ml��#�?�,�{y��H!{~]���x���������m�hb32�r�~���m���3w������\�����������t�A����O?�.N�cL�H�[L�|�^�<��yc��y��� �������x�����~�^��ˮ,{�Z��|0u�6�7�[�ٍ/k��� <6mH���`��am>:���r���}�6��Z���=�Ei�����|�H�i��lx�������� �����)8� �����f����[� ��յc����}oqzɸ�5��:�#S�YZf9X�)��km�I�����O+��Y$����@ �������Cɝ,�u!�����[�;i���q/����	N�
<�ڣ�U̗�54�	�m��|N�3IL�?��\���f���i�M�F�q����ļ�3�:Td����3��`��]� i����C*�ʋ-,��Iү
0_��؈��J�h��a�w-���ve�w����+u�m�o��91,�_�8!w9��m��v���[c��!�aJ�_:�ۡ��=�0���-Me5*���$���Z�O<ј[*�2��r$T���b*85uNA5f��{,�2)��f�t����U:�r��*zX��Y�����6�&S�+��G��.f]ɾ�\~+c�K��l���٤i�iv���u��ɧ���!�Gm|I����-��v�|��]���C�.Wl��~�m~��� ~	}������}ͮu��{��c�n���� �a���X�t�>Xn�/��>��[+߹��{[^� -q�~C���b6D��+ eѹmk������þ�ٝ��m��q��{�����`�~�����o��͐9�m{���[��~o���ؽ�~�|~w��Z׾�����:߷�lX�f�w��°�Uqm���~/o��|4�<�˛�2䲞�C�� JC��実e���T.�ˢ�6>g�z�bd��^��oo<S�]RA��W�c�^[M������(1��<�wkʲ(��	3�*H�J�z7�T�ç�t� #)66=B�\x�����lX�??f(e'�S�G�E�k[�c�k�s�#1�`/�.u�� �� LL��h���m�͏Q����(0�����$�u>ckn}ӷ}0�[!e�k}�K�Ԏ���5YCJ��G�q�$KΪe�Q&gu��ٖ��o�Qy��33\��D�2�b4#� I�ΒH��q�!L�+.�o���nT���M��>����s�lE���H�Ĝ��*�������mf� �X��M��"����LY&1_~����=�!�6t���K$3ey�*��R���,	�����q>'��&�H9bOBln^�KeU9֨�cQ	�)U��3�4n��X���1EYN=y�Uȗ��đS�cUV(�0��W5ٝ��8�>�,q�?x�5hL���g�lYrKk�q�oՅF���<�H�h
6�k��:E�o|R0a�S�%B-��$�� ��%U�u�ٰ��ǒ%�kɛ����>8��.l�`�R#f!%�`@kw8�m��nfal�����l��|0A6������2륎m;���o��pH����׻_���4%����:a��ݏK�Q�"��ݰX�l�mmu#_,������ \���[o��o��`m���}��r�ʠ[�b�X��ن�s������^�پ���ݼ|� ;��w�L\�߷�E��Θv�X:���q�oͰ;~|�k��}��l���s����2��F���ف�a��]��>@�������b�?Z�Lkis�߶;<j?;���{��}��{�fʬnAV^�?J� ,qa`n^ý:��ž���F��MUs�F�$�4q��*]�KuY�ٔ��N[��a!6�c�����T[!��1�O������ ?�b[���[���� �lD�������x|qU}�W��z��a�ya�{��2�lJۧS�[y$k�X��ms`;�������{����UY&i�F�{��)U1����l�G�Sq�R�o�$AGIW5�v0���7`�)���'Y@Z��o{.���v:�n%M^���� ��"8Bd+� i3G��SA=54�<	͑�7&E�L�eV�}�pF�s�d~������_�k�O�MKW,�������X�c��S��AD�4yN���_��ܶ��M�M���|08��?�|L�,�L�>Ox����e�.FmTe��kI(�9�ju�}>��')��<�B��M�k�ȣ!�'^�L��]f"��˛ݽ�3x�H��r��e��9�����/}~:1G[$! �y`��l��HT��X��vR�Q�e�zoW"��o���!E��ј1��:6[�����3����E�^E��E��{���EQ�Ǚ�#���{�q=%��"�7 �]���S��K�ۃF:�yE��!��mv���ۧ�}���|o�ȹ���o��Gr4�����b������[~99"�-���q�8�0�����l?k׿}��5�7_D�n��\���{۶]� �.-����?����~��nA���H�{���<��[y���|e~�?�ol~φ6��|�;_���0V���w�8Ԟ�m���Lu�m|~V��l�Q��~�f�ͨe�cqc�L|��A{|V�~��QfF7�'�_�+������"�\�rV�a�w[x�����*����ȭ�{�j�ټ���lC�5 2��������*+��3�E!\��K�a*�'V�+�ea�aه}�bNV"���<nm|aa�
=Ȓ� 0ʁ�$e*Q��2�de6`W����������+1�o��أ��'�4��ӿǶ*��Y�����[_ČW�c��xR䛰�������Ơ��Y� ��m{����HNY��>\�-�(�Z���\TTQ��#5(�t��$~l����q�9���š�f���XKqp�Ǧ���Cm��Y�pŒ�]s�#Kk�I朹�@��!���h�y)���FY�-�K&�e`�����R@a�����X=e��tS%�0[����'�E!ѸetQ��-eRTjWk��v�-
5ׇQ/o�M���'���4x�q�F#[<"�m6i�_᭰@ki� ����>������jV�;t��'��}�I]s\�*�W��iI-CQ�z�H�3�7,F$7ʠ���M.h8U"���d{��s�6�&B�9Kpo#�zf�<:t�� i�U+�QM<�m;ʬu�1����D
V0���X��Af:Z+�O��.���'�����=B�	����{��~�r�k����R+��X��.�s�5���S��� �q{�Ü� �UK�I�{����7J�����l6ckf �,7���8[�n.׹>?gق�)����_���{��9���a�uI?f/q�k�{��˪���w���}�A/�6�o,G��\��5��N�5����wP@'����c#J�����a��zRqk|�lx�8T���o�� �����{�-����	6=��������ϵט����b�|����`[v8�n6ǽacp7>^W���o����?��xW���i�`��|�����y4:_�톣�O��ਣ�5x�M3�ಗ��.��l~��K$���Sv������S����$� ��sd�T���Hx匐��U`E�!�A��5�P�&��:������*�*eQ-��Y��-�GH�t����x[l�<*�[G�=�0/� ��# 0,�2}�ܵН��#`FjI�v�u��f�M-� ���q*�,{r��B�j6{�o�lS�C#�"���TUr��n,|���/q���e�ݼo�6����}��@��O������P���oo�n���Z
�,1GL����\<p��VIa���{�⢑)x���y>Te\��M�ǵ�[X�4\5W�p���iy�D���ʛ�|��
v�����{~δ��n�����а?L��r�� jI�:��B���|�c��Qq����w��c�T�<R�7�{C�����b��G�j�0jIle��,m�,
��#��l{�`
1@�N�o� �#�b�=F���]'��EKKE.�dFu,�X�I%�zq�?�8��4U����M?:5�㕙�d<�u�@MB��!�^��}u���Ze��0!-�6|�*�� �N8�u�:�1��*xMtС��t��>�o
щJ+�k�ӄ�?2y�&I3)$�{������1��ږ�r5��x�b٤hHs\�@?[5�]7����el��S2��~g�����6��������p@�m3\x��m�
F�b����/s��k�����k�������������G���� ����[x؏,�)���u�����n��㍼��M�7��~��k����x���P\�om�}1e7{�vſF��	�y���A��.pO��������k�@$�`�|k�`��ck�?�/��� ����_��_\<p=�_��7��Nlͦ��{�����ًv��e�|6�~ v��]����_ݴ>g�$���fe�ӥo����]1���4�{:�9�<SG#!�A��a�>�=!������X��G+2�-�CtI�T܈�ffbć#�Ύ4*�Po�m��*�j颕'�.EuGd��Q�,w'K�=�� ��M��F�ɯ�B٬2'Hק.�~�߇�(�{��1�G�?�ړ� �^P�I45�-�X^V�s�9��R�H/��"�1)�D�4�`2��@'�(O���j8V�X�������+�W�7�׳dv �R檒����y�y�����n}�0�o�mqħ�`Ȕ�c��a�&\�mV��Z�J�c��S��RIy�+M�� �7~c]_�ٽ�i���ܛ�p=O+�<-6�v�;c���3��UP$j�F��v� �Վ׾\݈�*u��tM.V�4��)����lPDVK�GK�� E�X��{�X�KZ��n����f����������
�n�� ��������k8L�&�6FT��gO�R�T�f&���E�W��&�jUd�VY�8WVLϟ2�>�����U��Tը��3;G��
�u%Xe��t��&c+,p�ěd	��>��N�c��P�d���,���+71$Y@K7�|����xe�WSR�k�D��$����K���%���c|KOQ褼������r	-��e�yv6�f|���A�K<��j�6nB�$4 *��@<�c��2�O!-�^������h/�a��%ٶ�y_������\�[��/��k[��X�{x`gL�=Ơ���ndd_���;���_��x7�!���+��6�k�l�)µ�I�c� ���`��,���RvӸ�5��~|�ݛ]|~_v=��O>�á-p5;��o��:�y�.^���3۸w���pKh �?��#&�}����0#V��I�:>�a�{a�K����<>X���k�/�����=��� L��F�K�_M�O�]t�-�� l�i�>@��k��u}��l{^���Q߷bqէ��az�.�8m���ŷ>[w��A����q�ȧ/�w?n=�͘M�(؞��ҙ/� R�m���?�8#�!�ޕs��V����o?�����k�7�gM+^���C_-��㧺1�bU6
��˗\p���Q�an��@� ө?�o�= ������*�l����B�ɘ挭��D	؝o?_G�� Xԕ�Ĵ��n`fr幍��l���'\S���="� +P�cr��������lY-a����?,z�5_��r�R��ȶ}}�I�d^��H>��y��,}��G{�YJ-�c�]�Ǯ�1�زr�W%��F�#��{���Rp������$�E"�2�U>1�s��\TsKHb�W�Ϋ"��h~�Yi���O"mW(��MG�8;}3qhn�)�Z�� y<��p�Y@̠�HɶhϽo��ٻy�-g���*���f��ɔ�+������I�߯�==k�$�]]jo��������p`E���Լ:��e�5�EU@�s��T���}��Aƽ)�C;�p��ZU�me7eyn�vE���|��]��I�ĝOs�<����2�$vg�L���Ƣ�0{fH��@>Y��� ����~w¶m/�<����,�����:�`�b>W���� �������)���|>�,rU�2�90I3kbr�ME����51�5���!f@[$𾙢�)e$�/|:�����kq���X߷�6��uO�>���q�O��0O��s����������n�����?�o�O;�]��|����??��q}{o���V��;�1U6\�6��S���oc���q��pl@�S����[�c�7����[���F���2�_=�^x�Fv�v��pokxc/n�����m-��k��a��F�l8J�pN�f�T��> @��q�k�h7������ D_���q�:_��t��>�b��t��x������#o��6���{�,zI� �J�������P3�3'gO��{[���{��z4�q.	!���oe˝g@�Z7�nb�X��c�3��M,��9��MV���R7:�c`1ɦUe*�n���`um2�`	\/��TTdU��N�1Y��+��t�E��2�E��7�qJՐH������1A(�_P����í��QzY.r�J��O�ӧ���,Ch�F5]�e��Ð�<��-�*����,2	�Ji���L�����?;[�x�QT�Hx���+"��,��Y��a�Pmr0���!i#�g)#���M�{�s�;j��O��%��޹fPu�����j��\q~���%g:e� �=ͬ1�I(+�a�}�|�!yzW�P��kh3��aoc|� ���0N�lr�[l�H q���_�)�^	7�M�6ŻilQ��������B��sf*Yu�6���U�"Ӭ`B����FR�gϔJm�-�K.��~�_Ck)[.����%G�m�ndm|�����u�5��v#������MŬs�S���>}�ō����l�MΘ�醹�{X��_��a��'�>^L����1���0(UYY�d��^���໓m�������<�8����|>z��ذ(�po����^�~N
�r���~ol2��Kw���6��Ƨ�i���c��`��~_w�ǣ�#p���K�� +i��Gk�$�3������C��ı���=���8����ɰ�|�sr�����O�u��3ϣL�Ln�Sȅ�� �e�e���FSR�u���kx�p�9Z�VP{9G�:jk�a�Ǥ�� �:����~Ű�"��Դf���=Jw�x��"�-���2�p�'��&�W��f�Rupn"ܵ�AaK,�Z<���<�N�Lp֑TQ�QpjZ
�F:�$���8���u5�je��=�+�ʣ5UC:�Gy$������YB�@
��Ke�� �� >��W����3��T��ͮ׾[\�<��
e�gib�H�9�h�h�lH��7����ա6�����u=��;� ����="����`��(\��ë��x⽎��^�ܣ��ֶ� B�>V��2�\���ǆ47�m�2�<��[H��K�?YI���Ly���b�A�-�~��q����-��;��'� ik�~>>X*M��o��aË����c����׫��S��D�� �~��߾�i||�6�����w�]t��<����7�a��1φ�>���7���_���2*3�3_[m��ƒ�?�|�?�炾��|����y��?n;�|1|�x��������mo�����|�O�7ǣ�~��j�C�0�� �����<,1A5J�-%4�$�O2W�K� _\̬ŭ�*�
�>'é�	)�iK��đ��9��C���u���nV���a�}m�7�ؤ�Ҧ��� 2�8M�0O��o�Z� zM{�q*���!�V� sQ��D�('A{����mA���q�������i$�v�Pu�<W�Q�ͦH�m��8$�6fI��J�����q�?��ƊB�� �����a�jq�T����d?J��/�����vƿ�p��IW��PJ�_Sѡ��Ҩ�31夭0Sk���mF$ʖW2��`���[y�S���]�,ړ��]-�����8��?'~{` ,tͯq�
۔���;�2��>C��i��"�ų~|>�ָ�|\���E��5�l�����B|<�mu�݇�-�6�ƽ�c@>[�c����:|�r~7�ԩ���~��A��?<X�ֽ�>8�����X��R����邾^v�~8 XYM�^�Q�ݏx8�˷�_ó<Z�&�:X�?n<�>m��� �{�#���(���4����|6� f,6=�|�U@�~��'O�]����cѵ��PH���S��O�4i��>�t������(y��<��FT{�|���MA
M��1 uJDL��V�Mn� \��K�=$NS������`A;f!������E�ȃ_� o�*mm��jM����E�� �u#��_� �ܽ�r�����qb5 ��6 �o�}�� \Fu����~=$��##SCI������'��(-� ��lf��u}����>~�˝"�?����3^@قB���otq�s	�v��9ex�e�^X�av8�++m��|�#lT�qE��x�\�)	R'���&p��I���j�� �DԜ>T��y�yL�8^Of�M�ƽ9�a�nt�FђL����a��� r�8���'w��CD�^ݢ��j}���9�����ֲ���5��ᑏP���V��>8��hB���#�}�~:�����t��{���߷�:w�O��~�[�(�mp9-~�~��k��u2����x`4-s��#�4��m�,��=v�,u������������_�5���c�vo�0�ql�G\��Wԝ���w'� �:m��|�ň�a�k��1����Xm����i�X^ݏ|y[�pM�������;�� �W=͘���X���_��l[�Ā��}-�����k��za�[e�����H����C��2���j��1�~����b�
�~&�v7��M�Ӿ��p�`@��	$(�D9���Px(#���T��d$}e,��r���O'OgH�L�� -���1�!����#O����K_@���퇚X�ԜD�M`܉yN��\�i#t�|نW���9LDl�j�6I�n�|?!�*56���}�q�ޘ��7��tl�R0^Q�3H�ot�H���op댥����l�i�_#�� -�a�%��&�Z�CD�Xe��s�I���3eKZ�O��B�sY�X��Rc��C���
����.y�=,��ݵLdR�]2��T�#-],l}R�9VI)���j�����t�E�k?�qVI-]]M���j#�����Q��w�^������
�Zٖ����E�E����t��&�D�č�Y�����F��ļF�F�\,�$���X�fK�UU:���ҺD�b��5�zY2�+� y¬�ǿ����kr�93�$���������ţ��q�è�����#����co����\e�6b��_�u8���_me�t�@�5�a���s?�� y��a~6��R��l�I[���R�y_W��f,,��:���s��n��$��bF�0*m��}ǎ5�'_��?����Uܛ�o�>q��V��9�#6!}��هm�>�j�����<h��x_M>�c�{e\�H�%��� |o�}ر�#����0�}m�����[��<u��o���o����o�­����>�1��v�n�]�=� ?~-� _E�熾�����a����a��l��O��>����������0����\z8�eY#�asy���m��<^��W� /�N� �������lt����I���RF���5sS�X&E�r�:�.��*�:�%�q�]���ѐ<$t�3�2��ؙ�˒�T����w�8^m����)�H����z�}����!�J�ɪ)��i�ie��Zthr��̄��,/?�jJ�Jr��SH�$H�s�ȩuW��L�3^�0�ߟ��ĬNX��7|���������h��B�P3Z2۵��S�F�8����~GL��hU��^r�7~fF��Q]Z�j���E�&
�ť�5FW
�C\\����:S�"+4lM� 7	�Jd�l��en�Vp�u�?=��G��I9�V�0e�uUp[��^u8�b�(����F��{�Dw� �ow‌��8�r�����Y� k!N�����z�t�ձC��!���5�}.×|�@����� \�4Ԃ����a�J8<SVM��ٖ5BGO1��8<"zDgyNj��&�]L��Ir����i����݄��I<z��\G!l��;���G#��<<�I�Z��$�u�ćK�c�7Y�������zE��h��٣����"��⪫�h��Y���E>L�(�H�p3��i�'�i�]
h����^�V���7���ֵ�ي�hr��ƸY�5L�r�Ap	���a�����yk|[�8���Æ!�������7���?n	;�7>V��X�鍔���߾�����-���vf;}o�3(�O�Տ��N��;�c��?�XȤ���v��5�_����� n.49J�P����k`f&������q��~v�[[�a�s�m�le��׵��_[��kb��}Ʀ��K`u0���L8˟�A�}�Ǹ<'L|�?,f	��*ol]@n��:���� ,PYt~F3dM��6�K��X`�}�Ѿ� v����Ǐ�_���9�ru�}z�>Xm2���~{^�b��� <k�q�-�G���~�?D����Ǣ(>�=e�|%������lP��cZ����N��[�aOY��u�@[�\�ot�l0�;G$I�~`,κ���Ǥ�F/$�<J�9<Ѡ�
�+�4�2,o!u?O����\ieZ���cZ���Z�Hu�zJ��(�9�]��i{�O���$������AL���� +������� �Q��_�	��:�!�zWT��͔3t\�U]�kk���Z�wk[0�[w�m�QҴ�d��&a�j���,4��:⚓�@%���AF�,pb2y�-�$fɝ$k ��~_\���Z�J6I̜��.]���k��:~t45+�++��9���u��	0���������Wj�
���C"Ny����c\�v�9AUJj�r���}7�[��� m�mt����c�1�o�u�+��I�rq6��B��3���P���D�<>���$�A/��Ջi$��fNg+��$�]l "ղz��z=U"�����ut�㵲��kء�� �u�-M<S�Qq��lDrTz��\�P.�3;9������&SM<c3E6U�h��9��@�ۧ�������� DY��^E:��E���7�8��O,�:�(��WT��"���"��K�Ľ��+xu=HCʟ�QOe�k�kHr��va����Y���x$aי���-��'�����|qS�4T�K�э����0�0p�?�6��Ĳ�s-��i���q��k�q�|i�f���,X���k���4��[-���/���㰽��� -�x^������0��������li�������>�w�m5��^����w���R,Ys(�G��L.�g�����ƿ�������e����`k�<z��k�8*�2��{k�:�o��4�,]??w|e�N� q��㏿0#S���9��:�{����ƀ|m����m� ;��x��ë8nOյq!�6ϣ�걓�d]Y�-��t���~)�ҵ餆(����l���Y�3�e\�V6���������P���˕�ҭ��H���Q�)V9��)�4v�l�U��Z�E�˲��X�UAK	�<�fT|����cul�#�8�_�RSȀ�\H�Sv��"�I*�Q sv��G����G����,\�j����uY=���.d��6��$꬧M�]������d[z���0�UB� �C���lS�r<�E%L�Ώ]T���zlo�7�~#Bj�*FIe�,3F�#�e&�3��r�K��O�ʞFS�#	������6:zB2�����z�ʘ&��� d����z����9WNa7��.k]�huM4&c������q��=S���lu�����ۆJ�� �k�.��.Zj�THf�:��q�|��]��z���x%ON9ʎ9��D`���A��c�07ĲI�ƒ�p��S�H��<�a3d�	��X�FVճ�N�O:p��
XeX,5����L��Ǚ��|�/��L���Ԫ�ըVB�${DU$��pE����Α�M-<�#�𸪃��Ch���2���ı$kAYB$�Q�U�ex��^����օAZi�C2��wsu(m�5Fu[*�l��Oi/�\$��hc[�j[v#����DhÇ�e�}�\|���0:x����M�����A >��<�B� �����$��B�n�J�B.5��S�M�S�����yi����½��2e]G����=Ǘ�������¯���Kܛ|Fk1������Q��:��"�N�����Oñ�߃�K� v�A[��\7f���/q�Y[{�7��oШ��/��)����8���|hoc�����c����N�ƸSl\M����`���r@���`n�h~x��k��<�rn�|p/�#Ek���ط��������_�z��|k����I#S���#����o������m���_u��Ђ>'<����~�!�zI���_�Rp�H!�ON��|�L>��r�k� /_.Og�T��%��&Z�傦)D�9�Z�I�!�R��9걅����Zv����{�c|���'k�����*z�B$g�Guq�����UP	6�"��::C�ZX+��H���,���BG���-�2X��#D_���Q{D�V���׿�g�lM�\���T�BR�"�3��zN���� b�@�ql�\6�LUc�.Ge[��FO�z�]�������G�{�3S�� *�C��k�¢��Q�=�|l-i�Z��CĚ�F?w˨��|���5:�~�puڞxႵҞY%\�G��9_d��:�ݲ�8T�����'��/�9�eH�w��`����8�^PCf�'-�)�_R��ɜ�3 /��8�)>Du��#D]F�vl�L���9��/����<�5@��$�2�FdH�
:�i��uU8��h��F1ӧ�Z�]��B�T\^��r��Jr���4a~�5� � b�<N���	�J���"�m;0Prvᓲ�I}<�#��Ҙ+e��]M���ź�y����Mug�����B�,q�l�g�"�ԕ(@���%W-�>�/0�o���>�c����?o�� <h33mk�5�`����|�����ƤߟΘbN��K܁��ml1� �}��3����Z�?�|0�0d�s�8F�K}PF�}�:�ّJ��pvӾ�}�Np̙�Ȼ[�	�,;j7�*g�O���z�G,�FR�Td,�����_E��X����M�W̥���� G�M��	��e66�ö6�<���Nrzu��5?<��/|y��j<u=�~��o���۫1�>8X��U�@m�v�k�ov�!�dv�궲������7����`���`���ů���� L[q�e����o��q��ʛCxi�s����Ff�S+G�r�������5t��;�	�=q)��E`}�����ʥC<�#�;�f$�{xm�::~�n� /��2̔\r�yQU�V�t����I��V�0DR]�8JMGGYz�o2A[r��ax\e�,�QdȠ x�(�NYNo%=��r��5�+� ��|�b�j���W�z�eD�kCf̷'F�lY2�k�X�p�A�u��GM���6�[��l$��:J�)͙M�����┳.cOn���[�����ު���$ƋF:c��\��7sӘ�|�&�=S�q>/���<q퓕�g\�3d$�l�!����.M£Ub�K��X�K�br��V�76���3�����(b<6޶5$��1����ǽo���������3�⏃��G���w�ιQ���L�:��؛�j~#A,Us)��UC��u�c��6�v�����EG �!��M�o�۷�,+(X�b�9טX)9Bf�7ٻ����(:�������#����{�ŝ}�~ͮf�9���30�?6EB�(;����
���ԉ=j��b5l��(�r���x�G1P2T��qvWu ][��ƴqƠ����ys����Y5�q����@y�����Mo�Y��N�je��j�����oՐ6���:�>�����k���id�� f���?L3�zl{��Kb�@��k�J�As�I��_Wh��/Y��0����e$����Y��{Z�h��c#��O��Mo��*�����ֵ�2�7��V�K��{ƌ-k��mv��ǅE'H��8�,��c��|��x�yp�����:�o����F	<H|Ar̊���к��n9�VCa�qF�j�E��+���!���Paxbl��8��^e�Rپ�^�D�A�]m�k��4�����}Duq�Ѧ�|<p3YC�� �~w�����No�4����_^�ͱ�د�;�&��̨��;w>[G4J�]H+g.��g]��n�� �~6m�Y(������������Dsh��Uo���ǲ�k�Ǥ�L�(,�M���˯��xX�H�L��l�܋�w�[�lu��FvR�\�X�Q� ���;i�k��q�u�����m1�t's����877���w�~~��lֶ�._�;|��||��q~ؑ�)y
����i�:�`�}�зk�-�^Ň�]�O�pKӞH�Mt)Ɍ-��|{���������u�A�[�Š���q�.l�2+b�@F�0ۘ��ڝ�6�h�&���	�5���wmN���ƌ��M�<Ͷ��{bʓH����R��*=!���+��{HT�f�X}��6Q��à��8�#s�xd�c��߄"���&F�
�t�u�E�>-'
r~����='m�����ky~�
o�08��=S��jZ��5��e��*�)�ݭ��z�RK<�S�T^����9�����qYGW��
�/:��
��� �Kt��}̤��b�׶⾄|�,/�����4oI#�ܭ�]���~��n_�=��YR)���0[��\{.#�|�c�\"ݾ�s�w���׫���/V�����{v#Lsc➘���e��T�g��}Lu�Ž2�}����b|r���yw�� ��lm�n'��������禗?H�[�>����M�o�˂\m�� gt۶	n?��1���ӂ���Z�������_L\�cĸH?�8
����-�8�6��n �_����"�~����� O��,�_�''r�K�� . 1� �_L���O�i�}�?�~�� ��� �sO����\��ߵǣ�O�� ���,-e�\���l !@޿_���`��8�����#�ſ[�i� �>� �������?��pm>��� <[���K�G������� �2��ɵ�ۉ���ȟ�?���+�� L�F�B�o����=4C��e�|6�����;c3q�MK�Ǌp{�� �}���� �zcտ�_��7��ſ[zab�m��i�������.8���>��.��� ������{mĸOO��߾k�[�����k���o� �ֿ��^/骰������  �� J�:xǦ�����~����2q�L���ѿX�\�A���� �*zA靵:�ڒIc��㩾Oמ�1E+f��V{�[�oG�r=�slݻa�yx��F��><F@:d�(�E1|�^�"�ؑ���EjqJC!jw�WS��/2#;����h/a�'���f�$.O$��"�2I��	�F%���+�i�9��o�����7�??�� >_�E������H��m�ڭ�7Ƹ�~��ֶ2�7�c���v�l��8�o�um[%�9l�[���	0n���� j���!�]YO�bHj8�Sĩ(�)ᙸ�h)�Id�S���u"��:�/�_�ݿt޳�l�����{���=�q�ݹl�`(�`�K�EJ���� �>ĝ3
����G�65���/�#�Io+sa�������uzX�+��V�����%���Sc�?WW!>"�\�}� p3zQ�
�#��x�z|OlG3�U�<�+�*�$� ��$�4g���[�������l8�_����������m=_NQ+&Z���,�.˛!�̤i�_��N���*�N[)Z�m��H�(W�9:�`�F�c�!���rg�I���}zt����������(w�I��ca�W�N�YX�j��$�(��.aIn�s#H��j5�S���,� b�:kkf�i�|1g�E������a �����7NQ{�Ὦ-������u�^8Q�_��߃��7<Y������5���tk-�#��np��4�ݬsxaN�0r��P�|����-ي^]����l���.b�U�*���^��i�ݛ�pb�ĞNI����4PEQ��Mȇ�V|�e����k줏�i�Hb*#Sa�Ί4Hq-uzQg���7Ӻ��Bfk� ݴ8��<���^M�}M�I�v�^m���Yj���L�u�l�[]H�"�Q&U��1�P,HL����O�	��`o��4c[�>a���<�`$��[��oVe��"�A{��5��ҟ�C0��H���bZ��dK;�P��cUL~��Q0��dhc�����?��`���R�����X�%�W-��oTHPI�`�ն]գ`A�:� ��g���	ZM��ׅ�=�nj��|�d��$�V�-n��ݣ����H:b�$�
���e>Оn����A�3��ǣ�+3�<�D����:
t��1�m/� ��� )   !1 AQaq��������� 0P��  ?!��Ȗ��`�8�<Y;a�Ѐ����m���0����!��#L���*8z3EP$�C,��R����M?�H*��坦��@��4�1`Jp�� {@�iq���լ����>Z!,� A��)��_B�("��D�`�R�B�xM �A�+0T��pY106�T-p�����LL9�p�W����4R����kVb��h9��v\@�.���4�za� mJy4���9�5�gEh^��`�����4�B	|� �VW�*됒�Z��.���z
�&�y����sY��MJK1��6�	 ���ᛞj�)I���E��mKV.V�q���.hu�D��� �_�TA�^�M:Y��r=��$�P��a˱�.�ҋ"�"R��+"��b�oF�Q����8X��
�,�+�Rc��0R�x�	��_�JU\3D� <�Q(�laA�Z�"�D	_)�"���r
t�[i� �_L�1O�lM��.G��f :���
"�RHQ����o��w�9���Q(1$)܂J΃v�|�l�8D�UGpj��^Ru�bd�J
�z;Ϸ�: u��@'H��%;D�ps�yq1)�a}�R���}�8Y3�V��iÄӲz�e�yc؟:,��T���/)U�'6#	x�T��	��Uʁ�ں��F���0��p@*��V�U��Y�x�!��@a�c�8�R�IO�q�@����^e��R��
�'a`�3;(	7��Ê �
Vd�F�R�m3�	�@�t�� A�<<ܵT�1�h��[��B;	"�iUR�,��v��E�G(N�m::�ȥF x���3�Ҭp� �F�T8�
�Hrx���zS0�����H��0��煓�� ��$Y�������,l�eM����^ ��n~+h�9��sn��t�8W؃AG E V,�c�Ĝ[J�d��9rۑ|\	 �_G�����f���ᡕu��)];o3�8�P�E �?�8E��^�ヂ-g=r��5Ӆ��q�y��e�`�����Ԧ]pUCZk ����s8C�q���.8��"��*^�:(�#67P���X�a�t$��� �x�ڍXB a����,ZP(�C��;�+"j��G>KԒ�81��.�Y�����?�W��Y�U/.�Bf-̂1Ls-A�R�dW���D$vGL2o��zb��yAT!~I�ܗ&��JA��8v��"� QU���Wd��;'C�[��A��"X9��&*���A�cR�b��z�O�7���`��m���� `�����a�2 ̱0P$�9�S)������Fib���j.$�� M��t߰����źa0��H��!s�^'I T�##ۉA�C)�h��m�r� �"��X�DNp��\�PY���-�h�B����f��N�Jʮ :Q�J�2�,�B<}���Q�F������1#Q1���f0\k+(p`Qf�뀕�fj|�N��ܯ1k��a�ǣ�h�((Ә4�jC�J'a��IC4�^�I�G�Z�]�:0�C�`#a)I��"q[F�J�V��^��k<5W�K�.dR���dV�ۂ���I��A���d�~��Qr,�[g��8c�,Uj�� �����W�vl����0���\���H�m���	B��=�3|����F&|�t�Z�:Y�8Ġ"O �!���Ȓ$M�Q�+a\�p���e��f*`wN>1��C��)��<���3$��B[q�V�S�8�=g�v(�#�%j%�@`�Ԍ,�5�"z�S���v�F8� 5��B+�%�����5��r�H�Y+�uK*|ˀa��k��$�]��� nRE��&���A� #l@/I*jG�_\�6��w�e��2\¡	a��BS�0�T k)K���#2�L�H�-=�)�4h���U��)3�cq���^F���5HE���d�S���+\��w��&2�b$t��L�)�V5ڷ�C���"��L���� �]�������F�戴5
	́�TC�~x;����1��u�P�e��f��>��n����"up@S�S��zHҠ����W�o�T�W���0�P��1@]ųjS���L�fj�V���5�$�$l>����U���C�@���ɔd82���h��F�2�i��1q���̀�,L	�R`�l�#�\�]Ȉ� �)*D�*H��Rq�X��=�$C_6��Mk[�`�����������/���j/�vʚtʠ� �l`)�8gf���/���Q��� hj����p�R��6k��,hiQ�Yy�)�ѥ�:f�qn�%L$�
���p�� �L�ǀ�N��.N3\_���������k�H��Q/{Q��1�&R�E��))��Hg8�г~/q���n`>4��$:�JZ��y-s��Y�;�A�1OJe��|���`-{��U���D�؞!)c�PG�,�i�^7mw��%:�����@-� ���� 9�z��K��� �
�	H|݁\�L�f�Q9�l�qL�k�/kf|y�M)��$�`��=�v�� ��=�w	���}�-Q��>Ë�QA����k�;�#����㑵� :<�?���%��v�A�����q�2Ĕ*��tĐ;ZxQ +9/�U�ԓ��')�@)��
]DP�`hVUN,�Pٳ����Q�����s��Y`�pе��n8.|��O��Lf�r��趄��f�1� ��*���)y�ت�Rq"�x" �u�9L=ކ�M����Gy��f4xѫ{��5��za,T��pU�qL�S�F&�>�*�f����� ��s`���4% ��]p�,�F*�÷\��$>�xw�\��_�\���?�	y�� oNnxBN�S��B��%0�X�����!Xq�y�����F���N��!9�!����.�o���������P&eah�Tv�`@$��wk�� �i�s�2���ۋ�z�(�9*6$���&���Jx����<�f$��Y7����B�y��^&�G������+}l9+�Ptf$""�F'����R��y��]DS���s�r����(E3\��/Й�%\i��(
$�ҡ���J©�d�!�d`<c.qbY\'!�#�/L�����iiG��Y���{�;�/\��������̚Xa`qN�^[���F��f�3�KR Ȁ@�_�ʂ����3�`�"@6�Yq����)��1�a�������   i6���d�8�(lHY����Y*�Z8 ����A��lX7.8���3��'6J,�D� J�0��Ɏ�ya҇_�].N�uQ@�M.fX�8�<��ᩢ�r[�M��/a��{8�#�ƀ2fuG�T{�'׌�(	y`�c�,Q(R�!Q��z��8[�~S� ��E��눮0�߯��p�Yno��/FAy����'�N����bWy�ڦ��8�x��*<�i"@9X	6h�ʘ/@�)�����v�U�ɐ.XG	<���)�6��b�:U61�6 �	��0'3��Q��
Ӥf&��6� �f��s�}uv�z�T�!� �QW�������	F�ø�5��)�Jf���$��Q��:��QrWH�pdT$�o�!�i� �fe�'��/�,�8h8����A��uY�n^H��}�.���84oI��^%Q��;Z����!p��ʩP�%rcRx���M`�&���3����ci�w��,��Hgi�!��� 8�5si7MD�A�ݲ�c����z\� %�R^�j�V�ك鉄�����$哷I�7�p���S����O���$��_[���4~��yWk�����JO��m2�iǈ(z������]�� ��B,B@���+zy����5�C�@��/��?�7�K�y`M��\�o��*���ŧ"RK'�u�L��j�-pד=w��L+�Q"����0�2E{cL8�´8��N� p�K�0DS@�
O!�5VK�L���� �������E8��΄rd���T��r�H�) ��FgɞDј(]"�v��d�ș'��+� y)����Xz柒p�1��ׄ�
�Ħ��]���@A��]��fqKT�#��=�*#`Ix�E%!��Ñ� �,�
s]�L� /3#Q�3L�[me���
�K��ɚׄ)OA�*Y~?�3|��n�L�����[=�bs�2"�-����3և+�̅:xB�6X�6��
;ڕ�"�Iu�g>����`��1�&�NHd[	����I�-�X�a�$��t-:~e\�`Y,%-K�������)�>'H�%�T����<�!��8>���FԀ`-��>�U�G&,W]����,W W-��%AF��%�pA�$���r�$�r�Mu<���Ȝ�g�7��x5����eD�M����'�����1���H+� ��_*�B@���9>��agN�F�{ �.̈́k��x�fm  ��>W),H$8���8�R��f;���
�-�8 lp�Qf�����TU"^�F��a]���<�v��c�P��P����f;x���f��fxkRc�}�B�نѹ���<[�(䣃�+�d��8��Cru�{��(8�-�˛�@����-r� ;��b�0��M��$� ���B&�WX��3`H��B��� ��9�U�!Z�(QL�!��������z��^�К�,�7�$XG8y *�<\�jQN/M9o�FB\/�E�(����� �&�X<
��In�&�ea-S���.�7�ӖwSRN�)� �`@�Ŗfj>BE��NŌ2��hz�9mh yr+�pŃ��w��0�[P
��'���\t{>&5�$8��f-����yY�H����}d��Q��G�?���V��;��`t�
���n%"@
G2r����O{�ӧ���x�N�D;�Z�D��I�T���+T�H٧د��y��dW"��˄�)2��PmZ�@:�T@t��Xʆ�@���甒�hp�7�߮��b�w���z� r�j@}dB�i�u#{�ӊ<�)i�A�QjF�J�N�}��rhY`B?o]�}t�e
񓋠uL����G Ц�Xb��c��ю�V���c#�͓&vg|�\lpk,�yf�ky`�1�#S���n��G"���`�R��T#�J(��t1G&��A`Ĝ���I(b�$;x/�Z̫����6�Crdl��ɩ�3x�2�9�����%EGO�喉6��a�)�R���� %J9������� 8�zT8�M_��5xh���G�a4��͹3����6��Ԡ{�J9�y� %� ��n����<W�ǝrK�-�:CgW��
��U��a�%�u^�>9`�bAEEQ�9�n-} |'Q�������'U��56aϬ�<qS;�@�0.��?4�l���x����_kg�p�2�R�)Q@��.��Yp8`�b�+�9��w=��w� ٮU��4�d�q9�0�7�����z�S���H�x-��3C��ltR��8y!P�@p ND�9d�9U�b�@���8D����4�,2
@�s�
��NK�y�`�g�� �gTޭ��&�L`��0��8��S�}��MF��G��2SE��YU�é�(�R#Er&�ct���G�_\\��S���7	�	Å�,.������?"� S��X�|�)[<����F�<�\�a��m�
�.��av:i�@
��WJ�1��`
�Nb����m3䓘�T`X�a�96	�^d�j���2�-,�:�
H���b;���%�U@�p#�F\�+Xz@�ʯ�Дa��v�_|0�7ʗ�����e@�"�b�=u��@�x��VA�zw�{!:�S�5�,�X��vNܫx��\�<�a�I�0��YL@�V����ºpS���.:�&!J`"���>�e�a�s'�^�|#ţʢ��׏��.=ܞ����˞�}�>��&���Ź�&w�`��������=�7v��0A��^c:9�c���:��}c�@x�������2n$�#��'0�Ԍ�Ε���D���"ag��������䒋��&%���v���B ��&�M� �Jj��p>�˺A��� �h�����_=^dB��	��'�/����6��T�\��E-�u����9X�M�X�\35&\花F����5b�ɰ�5+l�4�(u./#$�R��09�?S@�HGߨ-��q���/l ř ���2��E��Q���B)��t��h�q�F��퐂!�;ȰkZ(!�	�zg�u�V٦�R�zjjӳS�'�>���,�b�H7G��Pt�a�ϳ�,��^�a�UC�dpW��4,S�"���d��R%ʬe���X���kM�r7�Z༝��q(�As<��q&"u#y���e5>�u3'�g_hQ%Y�2	�����+P�G���gF8��{�D7�.�-E|ϐ+�V�4&��T�B@��*�4/	wh� �5
��&���ܐ)�oa d����`�s�%�x]�σ�i��>&��˺��!8&�sJ�P&����-#8Ƀ�s��b�
8O��o1������pSB�~���>� �<2�a��s�|�'���m�;0���V�O?��_�3�����ϰ��́�6�j�0)%Ո�+FXu
Ǵ���6D��4�����t0H:6-�/%���U˪�p�?�;���}b���%� (�v.2�X*�q�N!�:D J�$�a�݃
�&.����0l�y�HÎ�ƀ�K�О� t���Ş���='G3��F�N{<�i�/R羐܉JZXS����'�>�:����4UF!���9qyF�#�LbG X���.�L�PИ�$$��n0Pq�{X�+�c}��� ԡ���^!`:��[,\q�kr��;����9�I@ x��,�h-�n�9��v�Nܟ.��FX�T�Ȯ	��B��h�7������ѫ�Д	s.�˷qY�ex{���i�.O�	8�x�Y�����`X;AbHU!0�=	k������ @a�2�(�@�+(�4��	\��*��Q�/� Q�=����B
NҦ$���nH4Q�� Uq��[$X���T��"���02���/q� qX^�	�ה�A�&�KZ�OH%$���g����`T�f�yQ	��PB���6�O���WK���\7 �PJv���ád�߃��!����S'Yuv�����#QP�qŬv� ]���F!��oH%��Ϯ"�t\^	�a_���5�l�#b"�^M`���.qEkS�.�1�c��v���ǃ6��u��9Gq��� �)�๕h W$e��,MnM�Xe"Zs��#J��9���H���\ޠ���I��
vct���1��YMB(@��7�d�2��p1����R��\�!�����h�Ik�Lk��Ƅ,f#Jfi �p�s���>)2��ѽ
P*�cpi�A�!n|[hgx��Q3l&��3�$0���$�ł`��-'Q�����[N19�r�YG�X��<�~@�4 W�rh:����q�r�WMT�4g%HBm�B����Zr\�i��q-��3�pG9v=�z��p�G�Jeϓ�a�h��p�� �
���=�Bt��&qHh���Ξ�"�1�.b!�6�,;~E�`�棍��y� ٟ��.��VZ'`�wf)� n�����f-l	��y�L�c�"�B/FDH�N�!�*���,"���:5k�i����De�(`�R�>�MP�Y�D��X�s"x� �Y�!�\���K�=�C�zD$�R6���
�q0��g(����#�Ӧd,.il*HC�c�!�/�l��Gg*ތY}�)����Oh��C �Ap<̅=~>9�7%"�܀����+L�8CU��ƶ ��3C�$`���B�
]Q����UɔoA�&T2~?�X_�\cF����g�ʜ�!@��Zt\�v���7�ٳ�c�Z�qaQ? ?O����W�k  BC��'4dp�â�������w˭��S+��[��c^e''M��Z���W&�G�+�@@�W q��ю�̧�9����!Ո�|��{9���F�l���Sj�P���F��4	.��r��K߾;�����'j�P]Ѽq��`�'�7㆞	� e��|��B�@�Yq�F��G@�쒉wL�cpe����>�e�Ȍ�E�yE�+���5��A&�H�� '����;�_d�3a�(����JZjN�jDi�>*s�c5��kSQ��?6u�ǃ�yɚ1�Ͽ\� ]"N$4ڂ��G�p��o(�PDoK��(^݀F�dN�pu�t�4�����]U7fEAAG�z8O� �	?}�D.E8l_џ��\G��_�"�|e>X�|!a�)� LO ��NČ�HғJ���p�d�`腩0�~5P����q@1�����a���4r��܍T�����V5����S�8���
=!bUDx�lȭ;��?!e��#q=4�ȼK�E��Ԝ�вl��X�@E�1�>��qJ����qFXgUt�y�a@���,�h�"i�����a�	��)��r������,|���k� y�����;���h�N`�KzYɋ��"�(�d5�rҰ7g00v!�s�M�aW*�ؗ�4��e�?s��,2AF�XN\�H0�	(�.��9��5WJ��:����`M���-иF8AR����++�%s�o�|�-+�6�@�qӸ�D�5%���C�_�]yɟ��?��'�qxZ����}��-��B�|~q�#w��¼^��7�a��%�+C�g��DR/T���"����<�b<��Y�QG
*��s3�q$7$�F�Hk#͵``�,D�_`�	kϋ�SZ
r!cOiK�L�ƕ\�|�DY���tz9f�wgA��� \7�^���W�Dzݕ)�X�Z3!�p��Z�d}j[e�q����oG	�%�oV����Ă���<��{�_����nL�pPt91����~���|���-�� �)�Fq�����s�d��� m�q�8@�^���|��F����B绹4m�Xp��-Ȳ�-�����Dw��hVSy`iP����|�Ss����7����-����������!��B�ο�x��Z� ×��p���\fq�揟���� ��D}���]��p����
������MF��32�/�*o@��e��ƕ�~�����8xE˘��!1����<�:�\���=����J8���J�`��
N!�7�DXD$��1=)���3�&�\����|�3(&K�IA z	6�19���W� ��7���\[�s��㺓�����g��w�k�*���o��I!qDt6'G��4�s�V��lZ	�lȝvD������^�i��%�Ξ��ż�]�%:�z{J@�����x>�[Sظw��n��{�*d��E� �x�3��8�QF1�����1Ԓt�l�M�,$�a(s�.����K����{��cQ�@�Nj����H�ꥺ��SZ�q��S4M�����V��(��� 8��$�����?Jd4�@%�2wX]m�[�|�M�'Y�vrej��>�a PpQa�'�8�vN��H7�fl0d���X��+��V������f"aDC�`��)���(���F�	"V+\a��~��߂�W�B�[d��_����k��Yy����?��<� ;��|q������� 2�s��N��ǫ���W��� �2�˻����7�q�?4%����B�C�\�Nc�kM�Im��0 �XNRU`'o��� 6�����L�-xw
��✾$�.�(Ln,��vi���j���W!�A�4�� � 1���E��� ����e8�.`=�u��z{�4��w~���Ǯq�Fe�\���&�� 8'��Y��e2�����=Eth*��aB��M�������-6��bi��'�\J��2��sɘO�����D-�6K��Kʸ�߽0�,x�jTC"�2��d���L� :Y��3�C�!��\��1�B����s��F(�α�YC��98��F�^��e>�B�N,j���iџ�f�	�p!���cr�Plڧ�}���(�"�%'qMQ9��//�p҉P�H1�~�-
J'.)�ZZ�l*y�6�z��������b��i�l�o�������r�c�"�4�[�Db���ں�˃=Qm 0�0A�k���i�^�6�����jw֎-�����/a��}s[<����s�lE5����|{����]^� ����
_��?W�t$�k���?�T�!Fp��s�M�#�q'�r��� ��jjF�;X�A�|�q� ��{s��B�H�^���QƳ��,_���d�x��:�VN##���,�Qn����`��x.�L�+���x�]�)y_�p�5���ˠτ� �vW]$��j�����]��B(��y��)�j�r&�� z�1�0s��=��_�5�݋�A�� N�;�6�)uI���B��0��������I��e*ܼCx#�)+Aɟ�dy��*Q��rӊg�߭s>]�y������!Y���q�E�F�n��-'�af���_& ���� <r� ���+w_�����7,]�9
!�8\p` 9@.�J�*���22<�`�e��[�S T
5p1t~�yq�aey�?�48�~���ש��2U4A�.Q^E����M���@�ּ�W/u~#��gqhdj^�'�����.$E(�D喙��L�px$���rNA1�"�����߉���R�g^g�� ���.�� �͉�_?<_�}[���c;���~� ��;��|ɝ|[��� ����ȃ���C9-Z-��-b�,N���N<�R�Q�4�z�ZJ �)��>/�{�䣼T�5��fʹ�|5ƪ��o��:@)�����û���yJ�!71��׾`��������������7�� �4�	`B��3,��d�~
%�@G�J�o��v^�
64�����2?���3�a�Z�3�	���|���X�C��x�*�A��3�2X�&b�_gB���LE��Pt�%!]yZs�����MÜ'�r\c��Rx�9t"�VIǨ`d��!�z�]�8�� �]�]z���u _��@�$��i�O���4�D����s�N>�*Μ�Cy�%� 8Zk� �ɂDp�Ȁ-D3;�L��qP`OqAʼ�V�s��!��a��o�$�-]��� I����!(&ڄ�16��T��UD�����/e�6[b�1'}b��C˚'ڔp��]1�%4��9��&�����}�+�Ov�?ߞG|��x!����������ׇ��pi���������1��y�d������A����s:��7��\�=z�fn;�~���.�&� �@ �;޾w���� z��ƕ������Ҏ�s��r�
�Iʩ�;��t^��s��������d��p��tD@�\y��%��4�&�����h����˝!;li�c\����yFL��R�x� y�뻽pLE�x�84V&oz��Log^u�ͦY�B�� � ��vÞ`�<��8���k�% �t0qdx�W����A���#4q��!�ݠ�L�I͂��O��q$ۯ?;1�F�e�aԂ�ǈ' ��U��e~BȨ���Vz��=��r��(�����$����N:�f���h�h^����Z��5w�4뉩WF"�}�l�k���폁j�q��-�2����|p��Q2�����)).�R����Z%*�0|�r��CN]v\m�,��X�a	R���oG�!�s��R�w�W9	��<ɾ�nA< �A3���zf �PlȒ3��8@C���W��qK��~�$���\�'���>����M3����5&�a��� �X��%o��0��=����ɍ�f��^� ��d�T��E�7�?|'(5��W�F;�X�:�ϟ|��&�ű{u�����k�����<�Jy�w_|�f����ox�y��V��p���J9U���.S�`m<�[Z���M��Ä�!�g�,�s?�;D5�hm��A� e�*�G��ƁqI�e =��^�&�5��	�o�q�?_�;d� x��\p�S, N��<}�J�<��K�"�6.�H��5�)p��ǳ���c����  �B�k��nh��S0�����Ɔj�s;6�bsHB������Pg��(�3�cpU�c�<֜��S�[�@7h�r�y4DY�^V��������O�灘Fh#p�a�2�g�����D�Z�+�ϻ� g0�0���A�c�x�	k�0�@xv:)��US���;�xq���k��3*q�|�}��EWF	9y<h�{�c8=O�k�����`8:BH�%� ��Ja�fhe���F���c_�v[���d[Z@G������Z3�Z�H��LP�Q��z���\��I�B��̨�hJD�Q���o��^7��i��ࣥ�bqI��������g��c��  jA�.�&�p�u�ET���*|%yx)�K�Q��7�0��(EJ�Te0.�f[��\��V��� j��	�;m�*�>��F�x�REY�KDl��B�_i�|���<L���.>tw�H
H��3���
�CGp�44^*���9�6@h"\1�*C��3ި�"'���$��q�5qe�Yq(1(`x@|G�m�\�g'�	P(p��Y&�����w�`|�m����E-�^���we�~9��g��Lk_'��Vu>�k��8��Ͱ��\�q|��]��X%'JA�O����,%�
�<�n
 8��s0�u
&]��7���&�9�DQ"wiL,�"1�X��;.<s�5�f`�Q~���0ኽRႲ�<���u,׍M�i�!^�s&��*;��e3�2�̐{YS@�N����D��c$_p����T	�ypg�Q�#�*�,��L�8k��zX�_E�#��{�eD�
��Da�N� 8=���a �#�t��$M�y��R]C�mpM&� ���b6h�(�VL��z�70��9<�o�PQ[6��[7V�ـ~8�4��J͠����N���H�|�*�)-�DW��1M� �,G!��U��	�D���"�����#� �=��s)�&+&p��-'�jcLp �d������#�ц�*H1C0�:���d�ĄA�����К�l�xp<+�(M#c;� �Jv.�#��II�U9� �a��-S�"��(�Iǹ�H`�a����V"p0��/<-�_�� "��?㿮,B�:��	A�.$֘=��y�g%ъ$�CoS2���ʜ[Hh��XS$�V.#�ђ���  B&<p�
SJi�h�+x��c2R�q��<�.' �� @wy|�|t끙"��#�5P�W k廞;0U�($C��ũJi�SC��)�+3wQv7�N�XZ��2x���b#�hTy����#�.V��*���6��'(�xN_��(��ceȑ�$�cp����ƅ�K|l�P
 ��F<�ٸj�"bq\\P�L��#Rv�HX$��C,B$�"e�vEϔH��L��RD����P+nAt���#���;R�)M�:,⪰1B�tZA��4E�C��Ӄ@
�Vd�Q�1CR�$D���ja*���G#����]�R��o��Sx׀9��V<�hPq�	�-���. �(�Lr�&M"�C�1{����U!I�����ec��c&m�gcnYDUn�'��	+�����E�	�1�TL��쇠�� ��ib�`���f��D��,`X1Z2n��Ĩ9i8i�kr��
;����R�1�5��wQ�Q��9յ4Z�a����-��	<Z��pT�'Ӱ^�j�GC�#�VT:;���5��Up�Kr�2D�lЧ0�U�k�#AIV��K�Q!��aA�-n:�C+���������Uh���_8�nh�4�0�:� ~~���7���x�S��z�}5<�cžq�k�ת'"���"��S�����sߒAt3@�8 `&/��? � <���(�r|rm��š?�l�,DB�]Ic�T�W� ��K�!qD�2B)&A(�pK�"�&S��]7��]I|Ǘ��n
�)�������.�r�t�	R�( p)�o2�x��iY ��AzhD����e"[>B�\6��<&�:��S�u"���r�`��޽ئ*p$e%��	j��pCҙ������I�ԓ�Wv0K�������W�@�L��(O��B�v�Y�/�� ��R �G,�~���pp�kb�	Dƚe�kBp�0)x�&�݅�Y��u҉W B%��,�W+![2���
�I�d�(sb�rĈ��Q��i$�1��Y�AMqNS�<1%x���eX���é��>�f p�-Ѳ�� �K�)\0@T�-+8�YD�fP��R�9�AC������8tB�Ş��=���+�K��ꢌ\a
Z�i�L�\���&�����5B���a��R���,��p�_J�� [q6�WC���ljלE˥��ݬ�{{�)�w�;�'�މ7�Q NG��;N�0k܃L��͖� .@ѿ����r������?qN�v�-��, ���K����R�Q�c����c�0���\5����q��
��x�(���<��k.�����|�H��5���<}(�윓�WJTj��=c02�paa���#��J�'h�Ș��gA�$Z��)��g�!�l���H(�����A�wH���0�Nz5R\�Kq�	^!��:��,V�ϷT�P�E �ڎ3��w�œdD��5B��#�C2�+���� ��G�&p̅j���$ѵS �^]��f`.�R�.q�k�������<JV�)�*��ba��}�fE#��|:�7o�k}r����T�P�b��>!@��<qV�P`b#GB�kׂ`H�	��0�Zb��>c�i��gKA��9�ԌX$ɯQ	J03[8Ʃ5�4��H��DG0N�S�k��d�$16P����Dv��r�$�E��t�0�f;����00��^��u�0A��@��ƿ`�?�G��r|~����] �����qX�0�x|��G挦&*t�q��;��c7�Sb�
���ߊ�����g�oHR�2%0����
�BhW�]�R��[�94�X��9���p4�۠�Sj��4�fih*���-�9���Q87������D��^ Nh\��~0��d�-ܡ��NQ��z��d1y+2��IͮO��`�r�p�o�KVv��
���J*[�� ����T
� &`$��L������F�_0/\��� ޹�o�T� �{pu��Y*����W� ��!��Eq^�=hY�k�w�����}���P����E���c����TPW�p�:���1`a8v���Y�v;�@�ss��6��HWBp��3��H�Xu��I�'	��.�
����V��lV��������0�����+�^<BX��xׇF.�cBz�Ǜ��$���q��@�0���mq{880�č����l�y%P�|vd�|Х�Ā(V��e��@�pc�Jo=�O2�*,��0��a5�k�clX���x�������sY�BvfFP� ��Hʹ+z�e ��"����zhN���X3=�׮:3�U��92�$!;�9���#z�a��X�"ޱ�����ܽL��`G(˷�떈�]/�� �|2� �28���9j�&��y�U��z)ɛ��F2���/?|�!p*�T�|v���{0g��;7�)�߿|����u7���&��=��� :(	�gˮMc�#��G�!d � ��<���jk���$n��|7�_��r�����%����� �-p���
��=0�:9U�p���_��N@ʹ����R�p/���?�pp1���ˊ\J��44��*�%iگ��H���Ji�Qs�N�`�\���W�`�Hp�Oܑ�`�@x�@�g�H�܈�0��k]rK�{�
PBY�P�L��k"�QȒ$��EW��	9~�� �&p93��ͭ��<�Z���sW�����0qR��)���5G#A%tS�������<S�3�@*a*0���9��JlsEW5��g[nw���;��\�p�!��|j'PPʨ(�b��>! <�M�]Yo�,!�!]U��ؗ�|y�$nGhnf�8ἠ���(��C�U�WcQa�m�TM0&�V�8wD`���m�dр�:=�s�=�@ś�İ)�,>��Fl�����0B^ f4���垞
�
j�a�3@&����jt	pBP(W�����T�S��	�9Р��!�+�7�eK;fަ8r�00�S)��y���z��LE#sN��_�5�UM�̟��w�;�l�V`�n�m�D�
�ޑ�<�
���&�98Ǟ������	�G_4�ϙ�p��l��C��,����/�������9�:i��'��������,|w~����B�H[��6
<	��:�;3��9���?G��8�6>��|��>���и%�W��8L%���h�{�,�V"]�}C��2{�??D
�p�ǉ� 8�<���rB)E�>U��6�B�~|�XK2K��/�:� ��8<D5 ֮ܒ3���]��ʛl��mW	Ɯ��emX2��_��qq�?�y�!��s�q�����C�m�f`�	HxA�wk��~x������ݪ� >y"P�g��'/�Uh^�+�@��4(l���7��o�^�v�>��<Q�H0���8'��)4�~S���cf��k�A��������sxm�S�g���*����K�I�Uxe	��+�y8���r�>@�1�PC��V��'*V�P��,��z|%����&!��1e���(P��j��K��ĩxU��������!*�s��n�C�3��DY��L�ÆN��U�H�$~�8 �	�~�����;./�&#�F'�<�Q��:����L3��٪��Z.LEf�@�L�R0~�SS��_R	I�kW�ͱpn@8Ű�ѐ��i����yrInx��L���c����F��t��^?���Iӕ���p�Љ��3����y��	�zEQ�c>7gw�PŎBȗY�<돛�Dt��8��e� ﾹ��,��H�X��HqH����J�� ��K�O�U�@
��2%���DR(<{�h@_I�ͮ%�H(�$S}r�(SS��N%-|ſ\"�`z����X#cȓ�x���	6'^�|�p�s���8�8b�67�y��J���C p,d7@�0��^��A���"����/�h�t�(�k�%#j�%b�,@�#�n��o�7�����8}�ׯ�߾*�+C9��l^�n��Ϟ8�q��'����8in^Od}8#?��`��_���T]�=��E��c;��4VZ[ +�,�*�e��� ���5��䇳[<�f��%���2�C��h;�����>ʴ�4J"���&�`mH��-W�s!4��V�nV���+�4! ��|��-Z�0n7ӈ��0M�iO�\E4@j��l�lZ{5��_S�	PJ#�����/��?jYt�s�s�Uݻ�y��r��f6x���΢ɿ�㿃�G@qMi�a���FFuG�_��9\�gt�ha��C��q�7�z�0�*��;��dt�w_nb�$!�n�o�+�`�&���L�"��k��RSw��y����
��\��!H m�
���z��iYI�8�t&����#)�ͣ�����
��8�B��3@cg����ȹ�<)F�#��w��+�v��4���&��8h�˘��x���aγ��=o<��)��ⵯ��F���<^P��q3�����7�����+t&��c*@*$$�j}�.��~"��x��W֐h��zp5�YZܯ�G<m��D���q_��<���W�8\)�d�sׅ��5ɐ*FraP��(��w�_aN�*�{궰�&0\șr���*k�����K}k����/fxo���9I�#s�� |ɿǭu���Ֆ^��jvK)��ĸ`�D��e�ɷ�3`��;�If��tg~x�<n�"���d�K��� XvӍU�+�Rq��<�/�GB1��n�Y#�G���s���?��)�0%�R��U��HS"�\�5��*�fO]Ձ0�C�@,�gw\DXF��M��N+D� ,e��,��ZL�6
ߖ����d
|��]wƦ��Q�Ӯ�'��D�k� ڪ��u��N1J�C�}uͬX|�n�?�Rt#�߾t���Ȃ�D�;��$5ڻ5 �U"�����Mra�������l�'�pXP��r�Z-Y�����pGb����덀���6�<Z����r���p`O�$Ç�� I��hd�FP�BIP�pc��p�!�� ���@L�*�x�*`Ru6+4 �6�;�����Z�P����(���k��1ᄹ��:�6>��y�)o��V�C��&>�"�(`�\O�V��a�mi�|)��� �#C.-����B�������T��	'�^��צ8�j�0Z$��;㩒'(g��w�bD5 �i�q~P�zӘ� <rXf��}>���FN������%p�(��G;�ZPlJ�6e��QD���zbmb���z ]̸;a�8nL��� ׾-O������Y_(�;r�J�r�^/��A�z�3�h��c)����2�0'^2sTW�?��@s%�z�O0�ni�l0��h����� �ǎ&B�ʝ�ͪk��I-ڀEr
J�X���C��@�vo*����p�����r��bO�?�,r݁jpQ�P4j`�8�X���l�z�i��g�z�qV��w\�W���#)��9_<�Q��\⺭���g�;Wz�A�a��0{�E�L#C��r]��v����P�����+�Z��Y�M�D<ƌ�F-��S��r��r�z7~�8��x�}�|pVz"�bXia]q��8jSr�;���X!����p�όLp@a�<��e��R� bP6aɄ(h0Q��xi�t�����C+�w�e���4�%��A��o���6�0����Y8�˓�C��S�/"�s�0B��1�˨��j���:iNT!�g��X0���� W��?`�ǃ���Z���뗿�1\�.�d��'��/�̹��˙,�^%�A4�+��x� ��G�$�1?�8#�h�-�8���Z�W~;�D@ȴ���1��?��%R\���\<{D�p���i�â��_�µ)�Р��#��p
���6\���L�T5UA��S�
8���-V�
9L9G�(�:��x*|�6+�_�C�)�����e�LӉ~=\q�q����e0��2s���Έ1�&\s�R���A��,X籶��Nr�s���Fl� �TG2�q�,��e�1U��AU�N��+��H��`TX�7�\��$�#{� �����k��9�U���B�Psn>�K��Y�T�شFB��8R�s ����gY�(墡.,�P$��S>C�B���i�i����V����<��f̃�������=@�eC�@v�����z��к,����xgZk��G5XĂ��D��k��|I���0Ly��<�b�=3G����F0����X�C�;/&��:�wB��.q-"i����%`%WYO6x���zu�<�
���89>��[+������R+�$/^ԸfV
�Ƌ,i�g�T����h�z����<���g
��;��>��_+׻��]@<ۯ�7��eg8�� �
_K�}.�w���q&[����j<#{��kfb���"��8�����C�Hz����E|!r*UN���_h� {�.�'��(�)'�I�}ͯo��%�b���c�w��&�#?�!X.>6E1����S�N:�v�a�z�gpșM�2�"���j�3�%���tB%�f2�ʈ�L!	��(��b�Z��d�-��0����xF)�ʠ6.N@K"-Ď�U
㪂\�@�	�!*GwkI�pZ�����ŋ�,#�%����)-�쟕t�\:x�*��\�Ф��� xأAV�Y5�˄�zk�boC�{PYj�|>U��c0B�	�g	� ����)�'+�G4������"��!���4^���S�ŐZ9�T�廥�5��@���q|&3A��N��.����Y@���͔��x����nB��� �
븠c���<�+ L4��v1^���]�ˎ��	�sFUL8����$�f{5~�QpjtӉWw����%�t�`,*,�WJ�|�
qٔ���PGKHY"y�<kE�X��`���fvˑ�]��x��x3�ucߞ _�� �<iх�G�#�  �0�"#�7��%S:���YB� &x��[��q�́��;� =:�bL�ĭ \D���9��<�t{��͗��nmF%狳7稂�Ǚ��8+Fb�?�@Q�8ޓ�!���с&Q�g	(̛�#����P#���mG���aTk�dmZ��	,3����=�6c�i�v��'�|̚��I�)Ţ�{i�t�S��r��>߁����9��;��� gH��g�����;�*pJ��F_���;��p�47���Yg-�j���9{nHG�7��V�!�B�##Ţj&E=��ڻV�Y��Ø������ژ[���|�r��Z�m�0#��>!S�Q\p|Ll�u��sƹ�c-�8)�#�e��7�O��<<c����hYe1$J��.�.�%�H�W���o4eG^ �'�(�"`U�)��Ʊ�[�m�醗 �ւ��0���\�v��y06ݞ�%���pE) ����z�Q��]b���3n���D'L�ᥔ��t1�r���b�y%3k�o�Pňmn��&���1� 	P��*!C2"α���VQ��@r(�V�A�<��W18�@��:־������|��C�R�]�������a�]�c?��\"��
�2���{�	�ӷ>$v`c�$9
�2Jy��5 WE���������<u�O\�`=�&���3Ϗ�,+��]h0���${�Mh��0���zỸ3�94�Q1��|�Y��U&�����0�2��1�
�0}��P��r�K��Ɍ�r�Gíy�����y���fI��0 2&�&u>9��M��ۿ��`֦2l���_��O~�Z
�(�W#��h��:ҝO�������}}�,�;A�2BK�: ꛇ�u�����A��K���F�Rs�H@�<9W�����8����xr)���N�*� �9z8�4��	�(����I
l��,'P�4�I�����M���%�Sr��Cf]���� x������6�\_�R��JG0�M~��g�;�=�f�>0[�D�� 
	�{Z��*(L�Y	�(t�zP� ����D�Q�����#��4 lb�F�}�(J #���a�"�%�)٧��=KT`���_oACj�,-p2�7� �g'�� 3ɰ���;0�*a¿� �kH�F�.S������O|����r�6���	�mo���m���wq��|� \D][AK;F�[� �$b�1O�(8��y�-N3���~yH�P`K�4�t2<S<4wV�+�� �Գ�14~�y\(��:c�玧��L�3�8>y5S6�cs���i�� ��D҈��pƯ�_ԧ%T� ���Lw������_�OE�4���_��yj��͍�=��1�����-t��/w�,$w��+��Am�N  ���"_��8�H؄���g��h���=���dBA��C�%��0M��x��pk�(���i1�ȗNj]@i>�"��g��:�ɿٿ/� Y��q�}�ڊ��e�:`�& `�m۾6���t:�|� 1�| >׆	� Lw���x�q��z����o��� r��~<x���hS��6`��<,�c��>\��G���2rx��d�3#]�r=Wa|��	��n���>�'y���ʥ�����_���^lc����]no��a>�F��`�-O1��VT:��(�x{Ŗ($qN)��[[��2S�"�VP�F*sBJ�RZ^g�4���u��d�C��"�Vu�obi�:��qaR�Ƣ�����d���Y�9
sZ�}_	X��{KRLs�@+�|��M����4� g�x����|g�Į�����\��!ɍ�9N��w�;��#���{6�L���Djٲ6;vOA�"��	�G0���TX��6Q./�|�lXӳ�}pXY��w���ɛ����g�m)�  &���>8O	����.G���]f�:��y�|��:Z�uٟ�"��A	��%F%P�+>x֩�\��X��ؔ*���tI�#BN�˰�\��=]k�qυ9Kڟc�� ��`���}q��h>��3�_ff�_�n��G����l9?�%�3�qy�eM��:bz����Q�g3��oA���J��1�W/�TcC�I�JVW#?\� T�Y��أ�����5�K���dI�r�+(M�q]>MN�ɒb��w�s �+,0>)��?���!Ƣ���a��`���+L��}\6����῀�6|W����T�eb����DW�Y�n9�����	ٿ�����s����m��/盗Ď�A��bp�]1`�'r�3l:P[�x�	���s}�ݙz{� �S�7���`�FXC��^Q��
��:�.A5�x>uz��B����P��~�W/4�-�2����!��]��a�/|Vg^n�x1�t�_���~���fA$uG%Q퓓�a4F��WS�ְ\�{�`��������H��O\�>��A�!���G��
��d�U^D'N\�:�0?|s�#3���.��2 +&�����6/�|�J�1!O#�o�Zs1���汷�O�㖢4P�Y����Q��yc��1V�L�HxU�ݙ����A�5�!�̉��N��<|y�c��c��U-;CŚ*)�r~Xs���ڴ̰W�0 .�ͳ�?����9�!e�0f(� ��1"ӭ�`�Ƭ��#���k�o����"@��B�}xw��I�-��{d\��9e������`w�C��gX�3|-��� �&G ��s�*fl���v8$G��Aʬ.x2A�*��-!B�G3{���{� B��@�ÇBw���)+�8���u�����"��,��(#�E�n�^V����v�vA�T���#v4��[y�����@�UvL�:gpz�DiH��u\�)Q�
���t��8mh�����;  � b,�����c �b�qe��3ʫ�2��NCp�v���f��NAfQe\��֊!P�B�c��:�`� �\�>ϮA��W\O��2c癓'ǎ�7���n>8�������D����� T WD`e��a��Ct$����`x��T���_|7�+Z�@T�ylF[���f"{�|�ms0�אO�JRo]l�rfd�A���R����<��A�N�N���x:���8K]?��h_�^ �(8��̇C~K� yZ6ztc��|s����^��+mA�zq���r8\����A�M^��z=s�2��:�;��R�Z0M��8
H^Xh@Nwb �� ޹���b.�C���ѳS?�Dxs�����N��2W�[熇K��+/�O5:�� ���>e��������&��e�� �� �7	.FS����6�
|J������o�ٟC� �� ��&JpX�d\f����p#��p�A,2t�p,d<=}p W5�Vg���6����gqEÙ"�7�nO	Ɂp,M�|gD�s��� �_`/ǵ'�� 8Q`2�a2Wi̬@ua��� �а�Tw3o%8�����5�`�P�q2:���C�2�wys��PR�P�� -�&�~!�P��Ʌ���Y��+e"�<�M��us��T���?�GH������r0, T���<t��p�`��&)�^��s���W�
?�~��� ������|�����s���0*�gC՜�͊$�&N�\(�i#���޲�(�j�xrnM��+�"��5 �Q�a ���yF���2hR��u�(�T();"&��v'6W|�q��L�=� _�&'3��ʌX�E�8Z3 sF#'� ��Cj����$'��yX�pPB���);UE(��'�����~�g��NV����" ���y32�N#PR:9w��m!�yc��x�I����㘒��>|�F8b�㛀�� �y�|��
�o0�Z.G����+��9��3�a�Z�z/O .K��|#�c��� �8)-(�F�sxB��S����d��dω�xzai�9prD��`�����m��+^,q@|�۴O��"��S��o��	ҙu�٬W3�e�dn�ey_\<vG��J�`���C��<�Fr]�8���"s��u�-sg ��{+o�Y��@:4g�bۦ�x4��q<���fHc?����I���>s�tU2꯭L�%��5/G�'.��/EC��8Q�}Q��c�j#lGx����<�L�<\�`��^���)
��϶b�W�̳�[�|=u�i���~��HrXHx-n2GN}��.l���-�zXgu�l��ha+�A Lv��!�8��s�� �֩�eɍ�	ld)�7+x&`����p&�Q�Ѿо�5\I��W���h����� MS��T�&���xH2q��VU(:q�􂓝�AM*�WB���\O =�2���;g_,�f���&Op�csjh��3O�� x������]e�b(��W����A�Q� ���N�8�B �GB!�p͂i<�̣��״�!�����DTČ��PmEp��8�)�b֚Ԧ|�6�[2��o��W���H@ǎ��g�<��6ZC� ���!����y�4:{��ݱ�q8�v��>?)� �����_�w���3�Ʋҁ��?���te���m`�3i����@��;����\b�q!���g�<���w������)t��R_8�W��e��p`ćh�si��u�dR�S��I~��' % ��<�7�����Gd�i,��8�NИ��w�00��>����(y3Q�߾��|�#S9��VU�7ߧDUw�Y�80�|q���JLْ�'%������VT�
�}d�V;�0�H��%�+�:������0u�::��]�*
E�3R�qB�0��D(T}�8s�S���5��]p�����$���;\���}LI7Ñ�Y�R�tz8���.,�7.9w��2�t��4�����~-�������+���6�u�w�+8FjQ;�3�J:�f���Z熥 �Iw(J�� C�x�H�F��{���yv�w�u_{ǆlH���\J� :Y���x��.('2���V�q�{M�3~ �� �z�ʢ����Q�KǄ$c�`h� �|�s���\��ك��8��H�3�$��
il2�g'բc��[�w{�c(D��*�����y d|gϞ�$��Q�ˊ��8`*�3�2jJ	ٙA��Ŵ买��<��̀$���e��@`^�g �!�7�8�0r�t��|�8y":�>	]��;I�ZO��������e��� �Oɿ��瘐�!s� w�Ƞ�z�>83%ȏ�:�g���Ld2���E�mp}7']s@�o�o�xLl��N�.�g�Ƹ��!.*��f8��)��:;�>8B��Xfn�9�L��-��3�����Ǡc=��x/�,,P��&��,<���'�n�����w����f�$q?��Æ5�O~5�t|��m�\&�S��4IN@�E�cf�V�_@�j
��WnA��8�$��R X�p�a���r}�����=0��m��#S���r�P&L�5�>x;J�t¹vu<癊*�B�b�#
�K *���j�:ZC@j;׃���SŘ����z�3��x�����Q��D%�9x.Cd��"��*O� $�s�7���� ��O�2���\��Ɍ!H�Bθ��"� p����
M��Ofk�;�R�aC
������54|��ʗ�"�HB3��"��}�|�� �[�	�� �������9 / R�JFĂ38�T<H�fO��ʎ�����K��3�JK� 5 �l��DDL���a��ֺ�\��g����Z��E���*��X٘���"P���d�1�Q4[��Nv�l���/ � �x�.O�/�+�A����X�i�F�$�nc��JO��0��2�?�\����N+o�"�����5Ύ�����㊆*�� �y%�V��5�;ޛ���4)�V� �$��lDY�ˌd����� �l�a]9�z�!Q�#u��x�1T�@�)�7�v`�����8³{��b��"0p�i�M���n�$���dP9e��f����	,󡍐�vN$Pxܬ��� ��%������$~��:�YL/��g�?xS�,Y����7Bk���1��\�"?��mm���R�R�9����FP1�$�)년t<��.��+LqrHeb"tqo8 u��pC�6��i��*;	��\3"���� =,80`����ې�#�Y�ѨR��L��S�Dڌ�ȇFd<p�p��	��޿����h�wq�+�@5sЦ���q�tW����B�#$���*�J4pF�!�<q>��sK��N;�M. A���yG�PN�!�$6��Ff �F@�����r�M'Bʇ���+��կ�~�~5�������t�H�P��t~ ����l4��n,��<��9p*\fx���C�C�^#�o`>�'�W�V *C����,��_�3TV�O�=<S� |����8��Ü#�r�C�gF�x����~�X �.N\#��q��,�"�]�� �_�yB@���<^P� f}~-<7�6I�����?��	ҁ���8le� ���֧x7;��7J%��^g���r����9Aa��o	 v���Z�ĸ0�ί-����Y��_.y�c6$�D����s���a�}��d��u-�Q����qT2]���
o�y���	�֫��cgpXw��q�)��&Mjw���F����3#��r��;�$�x/k�.��qR�]7ŁJ��K�	�z�6.\8���#��zc�qW�F�5�5��ֻ�ֻ�Q��3����gD0_���E��7�>��bG!��`aSb?�~x�m��v�=q�ud� �X�As����BV��&�Qt��O��'!ˌ����o�))�o�����2����rf�PG�@�k�Xu3�4a��v����f��Hv��ǌNT�EL[�����8�:�*d�&����qQ���J�
�x�y��	�>*ZF��\-��H�T@J hf,ܕ�۝���f���x����7>� ��[ N�����y�Oǂ�l��VEڑ��0bP��Ts9��6�b��É�Zk8�p�u�N�L;뙌%��*�r6���(��/qw9�Q}rǑ��ً���%U��O��o`/�}<�����{�5��.�3l�^�Q�	��/`��V^ԫ1ߛ����vc%�^�34z��A� ���)��H�d�����F�i�ߊ�#��{�r�(S�WzyA
7�ju7Zq�n�A�|a+ �<��|���,����ĸ�2�sbz��d�o���<ꅌT�)����{T�jV-�L<�ES;gX�>8�6�K�C.��N%�H� Ώ�U�8fہяW�LEv2zCm��{?}�^�� �8z,e�\ d�%��댋 �y�j^�4���`L����lj�]FehA�9��ZJ`!�<w�Y1�l8-�C���**3����� ȅM��v�6,'��e������fE��z�c�Ïӝ�l���L����=��dߎY-SP�AP������5|�� *Cdņ4Y|��������L��?�f�q�1��/�5�*)5�u)H��)��Ev"�-���h�p�!#�J�&�: �&�����$"�-٨�s�#�T$\����:�\f������>�8"Tb\'Kb���,����i�ղ�eU�a#(�y�f!�W�����z?����������~U�A�L�j�E���NDqkW� ��2G�J�bT��T0�93EwL�"�:��F�s�� ����/A�R�[� c��M��j��8����#��E� �q��y�lE�5p�;�����tH�=�x-�'��� }p��a/,S8=r8��8�˞a#8��q��:e�Ў�0�8���N��T�}�:4�'����0��99��� /�	�;L�5g��o����U1��Hfd�c�s��쳁�����h��k��+1���er�#L���|ת�E+�i��<\�1��hha+}M<�)�*Pa�8�Fb��c�"�!�0����y��)K���@�țˀ���cq���J_#!��(X�B�V�T0D�҃��\ RY�k��g6�y\Y���M���nׂ�!���	6�.u�]�FK'�^�41�`jכ޽�ڸ|��Nʈ��� �����kqB�;Re��9�!:Jc3 L*hy�T�8&�+��a��.)�L����TM����y���RF�#��v�<�f$��h�bs�je0�̧I������v���B�MS�W�������&���k�
n���X,��y�(pl�`b��5�����Ol����"(H�US�&g?���<S����|�ldMg�s ��0�D���G�����q�1c@-�qlb��������6 �h���9+����0Q��R�U8�gQ���E�s�Ѽ����\2k�{Xx���灒"���n�^DS&D�2 =n�JXL.��Ř���u��u: ;� �')0����-=r�b���'Nx�0���W�� 	������WA(�&�$Ǯ6�3C��O^\1�#:E'����2��I�<q�A�-�[��� �����9f�u��ujä0��<��#�;�LO�~>�K5��>�<j]����)�s b�Suz��.o!��N���h �Ɏu�xz;}���\��`�?\��fQ��W���U4H�B4�f�c�z�p����4�! �q!  �\�k�����B!8� P��{�<��Q`���>;��+�g�
l	{g� ��v�ݵO:��� I�A{c����T�0�Jk��eA����;�}�jg��p�3�ק�7�ݦ02�dd��:I���_O\7� �
wLWyf�y�SjH4�M��02���9�5��qm�	��(/S�m�}pT��TO�l1�o"h Lѡ����ffq�}怼� G�w��'�����8�p�v�|c� ��!}� �G�
Rc7u�ZaLr0��x>�-���:߿?����j�Η�~������IBl"'!\�Y'�>$��.�{ft3���pp>B �-���`"1�x�g�t�x�+N x�Ο|��X��U=&:�A,�%s�VG��&��X���g��	����u����M&���(DJ̼�ֻ�>�-u�{�lLp�T��Jg: !�m��Q�88a4���7��1�S#L��3�� t-U7��|�k~���%�w��W��o�F
���ݞ���g�G��}���� ^,��.��-�`���}`9bB����X�� �)�����=q��1^��rg-|��?<D�9w��ߎV*d�O��Mx�Ƽ��p�p���L��Y5�"��p�k�N([ �ъ����R�ቕ��w��p��$m1��Bh$d��N`�+@R�ߞ�HtW8�f��"c>_�߾x���7�D��o��@�Q�x	"�:��B��Ƣ"%��S�_��6fv$ɳ9O�U��!���EB�%��f�\4X4En���*��:�
I�rV'r�V� �/�{>5��`
% �ݥ�)ITP�����pʏ��&'��d�:�6��~��oCx����� %J-�ɁH9�*�����@"��iO:�p=b���0��g0>��ᄘLÔ\�\0u)��6�����*�.��:�� �*^@"8�yڠ�4��*���20��0p��V�_[�a�Gg|�]��|�3��Hb�� ]��4�/+�:��X��,�KjC��NLp���a�`������Q+��~\��B(=��#�ai���^���Z���0���VY?
���(�D���������,�P�rE�P�֖���:6� F��5�rMu�þ���1&5���117�K���p���}�k<��Y�r�ǎV�y�kߧ��h�nLQ�w�:-��K$��K6To� Fc�`�+��Y�5�5�뎣y$��F����E��c�p��3��^3�lM<l�*�d�R�[<��e�b���r��:�>�����4�*gȾ�
�FŦ������?F'����1+�F�H!�όxk�h��5D�'�k�8J�2�:5.�����Oi�̜��U�%��_��|�t2�&��8A�Ǘ�x>��z���0B��{���*R4�w�ny8�i��}�(T�(.�q6j����M'�jq� |$�����	M��\PG)D�����EQ���9�_<, ���V�r�@�������� 5�pj�N	��>��`��W+�}�kt�t�0�+����B�z��:�8C�#t�J˔�l������xx���1!d.`C��6Z�A}���V�<��E��T�?,v�O,��
p@ �{3���x��~����o�R'䏫,��)��:5�8]@
�=/,�c���;{�ck%j	��&9/+Dn��dw1θ.h��v�N,�� %@ڿ0�a sȀ@شU�9�^�fUGQ�޼|DT��ޛ��͎��&]Pgm-ϵ�@�#1��⒏�ߎ;�M�n�8s�f��{�f�;��Q*#' �vw�N�B����|��x�f�8�����|��X��̊7�	r/��|��O.���X�]f���<,�g�9�>9�?���U�N��vz1<�<�іh���'���ƹ&�c�z�Q�T��Y#�/<��ͫ�(��8�W���W��Z:?3x0��u^�Z�������������!\>}�o�q�x��FX_=w�u�D:1���0%��D6�sO'����0�c��p�d��8i,9��_� �m�8�	�H�ݟ���|�� }�8f�τ��g���4����ʅù���w`���/	i�-F*�����A1��1�u�� \�� x��u���r�dȉ�C���0�5 #L:�g��:�%�'���6�6�1��R�@�6I(�00��n�8���0��D���<ă�&nZ��V�HzV1�:r�~2�c,�4^l�C�5W&" ڨ.���t� \���9t���th�����9�+���pO	�D37=	\��L��D�Z%T�RD5%rc��٨����y�[�ځjn4ظ^��^��~�x��e	���� 4	"x��&aw�$2�8ű!�X�/���қ߁�:���b�p��#���Y�4���� �x�"<cGa�\Qôo�@�� ��\OMe�e�x�7��N��Ǿuh�D(=��\. �S,E)�u�J �p����>)����b� C��:�R�� �y֫��ߺK� �����׎�r��De�9��o��Ꮿ]?9�|Ky�lY���n��� _�h��N��~�:�nmƸ!�?< �}7+�=z�(Х�`y�y����%��f�4'1f7)v��=sA+w�<�Ne�XՋ�?>1�s�!Ԛ�У6q�j���|��pOg�0\��Ѭ��ש��u'2D���L���g��7��%2�Ǳ��N�+��Ƿ�x-��o}�Z�$��brJL&�j# ��!���2�����3��~�4�h u���������P�0wگ�K���|d"�\:9��<��3��!�d�e�k�R]d�F*��z�������n�M�L�0K�n�X5��;B�yF�� �
) '�ۈ���8��!X�N�{�����H��Լ�$RT��0� 0f�e���H�{�?�=�����yL&�t��x�'��.f��+�s;�p�#�᠏{�.L�M��$���c�{{[�$��Q����C�� 8��@n�1^RRm2�C�.62�c��De�p�N��-��aY>]�sP���7ʷ-�M{0N�x�7�_��R8���M_d���y�	�3q�~O�����X�bx���r����|���38�t�a��$Ό��/���3�>�qz|�=��\2Ŋ��_�5�,��y�z㱣e�]��p�j'���g�����9q�69T��\p6?L�]��7lw�क़��;�|z���!j����m.<�?n`g1��y�B�	�dg��|nU�Z����0=�\���PXj����5J � �(�+��P�l-,�L���a��9Q XJ�|���KL�?���
['{�2x��>�|A�hC��TOPk �=��THP����n�x1��;�=�6<�}��ǃ|v����Z�{N:ZZ���Q0�uDO����P�)� ᱡve4���+ɪ5*}lB�0
Z��f������@PD4�ʡ��Cn$��&Ԃq,j퉂�!���b {��a&�u`&Ps�PD, ��8��p�|~?�| -��YOe���W���y�������e�fU#,A����lz��%ǎ>dJ����ݭ�|�{B��0v�"�y��ex��d��;f�����	#��~y`|��8�d]�-�_eQ�e�- A��O���JĦ�}i<g��&2�.h�ã\h�.l1�9��/��8�p�FZ��x2�t����G뙂��&�����B���u�}<�ʒd�2~L��(+�u��W������zA��|�D�B�4���s�/���	�ۂ��L�^����;%�-��^,b�������m�:�W��3�p�<y��o��\0V=��&�c8R�br�b��F�w�x�Q��~TOw�0�����b���ŽA[./xE9J���_^�xK�J�) 0������+��Z�c��.�TN�?�p;$�yͽ���Tg��3Md��`���1z.����c�g�冉!�)��&�IC�⊊�-�P6��`hƑˆ:��QՔ�1�!��mU4���Ȭ�P2����t�y45�������f���U����U����Qp���X-�~��?�	1c������@����<���0�0�i�|��l�  p3���s\����#�6�bM�R׳������p�Ka�,nA���o���$��a� !��w���S�??�t������}޸�[�.TX�E�7S1(Zo�f\A���H�\��s
y aT;��"���$�.xpa��E��e�ŋ�Z�'���&O����wA�I�_��SAp��6�>��Ć��N�}���t���~����	�����W�����9�Q{�d4F��
�W*�}��$��0w��^k'f`q��gBv)��n��w�k:���UI��ҙ.�
-
��)$�����)�ω留��n<xo�  `v�:�䡒q��
�T�fk���aA�N�y�t�u+��癗v;6M��F(���q�*��������3,=9�%r����gn�� �(P4�2� ��4[Q����M���P����^��5l� ��f��AB���¿�
f�(9�d��n ���� x��8��	-�ύ���S��9H���ț�)2�ƅ���Ɇ!�����>��P�o���0�`��v@�] � ����?��x�6 �ՁEu�V���?LHH�q���5��[�\��	�
��6wK?q�A����� Xlj��Q��?4	=��|;I.���R�H!RG�6�U�y���Q�i�b2i���\��LFG>c���x�c3����l� ���$��iAv��s�� D)��Ɵm�9���o�g�#�� �R��|������0�۸q�B#fbV��0�̦��(��;Ie(���}g(#�K��|<;(�vУyq����6'��S���f`���$�Zx�3�Y�w0�+4X�E:Iw�	z�z�8�����`��o�86b�~Y�׍[fLN�<��p1@Ǩ��'��XPĘ��+"��=�y�o����B�'Y~8�i�V��{��h�h�qy7oQ2LT�0ƞD�.P;�>���� ����J�&W}K%g҄�^�/p8@����2����8��~�u��ߎ�?��I�
���D�5��"H��5SD{-� ������� ��zSB{����(���t��pbtE�q�<ltv8ZE;Ro��}��]��|,ψe\��;�\H�3�1�
����yh7���~g����d�7|�+��h��[�.���}b%V�7m�P��v����d��fg��8'�W8D��6ٖ:L��0rF��*���\D�d������c���@6��u�z:s���#M��?��s�(�J�[�eHx̿>�H�7p��ԉP�����_kPa�T�#�!\a��ڣJn��bj�ݛoRFֱ��0ڠ�#�p���� �x9����^/��<=�!Q<�_޹mϟǏ���':ZW��x�>!]� ���N��'E�h
%=�	mz
#VS|�k:�ε��u��YlcK��.�� ��p��(['�ͩ��\�%R�������uy>�p��R�6��͠�k��#�\3�e�i��2���� +&�^�=9�a��DC�3��<�4h
�>x0����������\�W�k�^4�v��������[b�]R�f����,��� F�����`	4p���yNIA��.1�^,���ͮu�}(��x�j�T�¼h���˭0���!�� �D���^v:�G�7�Xg�z����ˌ<�2g|`��~��o
�)��ん����m����=�����	��ǖ�:8�Z]瑃��D�b0�2��'���r�e��ˉ|������p���,��R��-�S\u�Z{�ar/�`q�*e4�'�x��n���
��I�����7�d�;��	��hZ�Jx:�g[�J.7��(j-�"5��<8'$z�<�k#<�{M�?���?�^9n_����+�$���]�o�0��KW�����u�8���v�!*Â��LAВ��9��0��.t�9:�e?���Z����;�;"��T���S'Z�qA��,Hۋ�a�z�TAg�U�p����%�M=> ��C9N7�7,뽶 aq�u!)c�BX�Pl����b:�`,�7�b0�_���@⍌�I�<j��g)��~Șd�݌�><ped��q���j��22�?T��C��u���}XA/����.?�2Wy�Ĳ��`b�g�:�^��;�DLŁ�2�|�T�x]i�s����g�]���Ea�S4����3�Y�B��t2	����� ��2n�)2�޹&!rL�1�{�}�1f� #g�� ��臃~xJ���wn(p=�N��g��A��W��S"S&v�� �9,�+s[K8@ag�5\}��Y�ɝO�L��n�9�]c�<8m�3��֜SxǞ��(��o�xU(Fm_�9YĳJ܍��Y�;�fNߎ'�A� �{{��S�4lL����ʤ�&q��:��EP=�Aa�CȠ�g$ᖣ�QnY�m��e ����5�y�ɕ�3���ϓB��_f_�7`S(���\�{L�_�&��q�p���m9)�-}�P��ට�ĭ]AA��4nG0����8��/��)��H�@�4d0�(��$�c=�PU�u��Լ &�3BgA�/�ENH�*��O���9 *)��m|;a��gHM�`�)N�M��4 af�;�2:�����+*���,���WU�.�C[�"7��8�LQyJ�%ɩ��$��~X�H
xIH��(־g�ʂN�r��#.��B�P�7*1ZFTKE�M��f��R������/σ8�w�p�ڢ���z�S�H �Тůx�/q���< �.3���Z���� A���0�{��|��5�����+�یZ_]y�a0ݧN��?\�(�]����\�=Y�۳57oK��P$Z���"���%�N%�GT�55�cw���٭����o�p7� P����xɆ!�Z���`�O'��c�����y��<	x���2	��5�\0���[��81�9��D��h�(�=��s���(*����;�O��k���O���=�۞���[��� �Dޙ:�����cCE�͒�Uf��x��ψ�����	q��&'Jy��(��,X�ˋ,| $�U�w�V���וE]߬|�}k��������+�T�YK��m��p3u�C �<���@2���B���{�G��8�[!������w�/c�.q-^��~F<'�� R ������a�Eb��q�4a46)A8b��αaŘ�(緝k~ӵ�ԔD����'���I�]����'��! �(����Edf���A�|7s��i�񄞹���%����CEЙp'\�����`o(q7�S� �a�K�m(�j"�0>�>� ��.K�BT:���G��(`�@��O�)D<NEJ64���g���a�	s@"��ܬBr�N@�q2�Bf��df�ΐ����]i�Y��H2�ng���P�J�5�7��lfV�!��{q��\9o3' ���@�3�S�t*�-E��v��_9��	�#c�� ���f���M��N�َ@��u� ��ܯ_�=�\��Б�o�| TI?���m�~�hZ�fvx�ry� *�M�<�<�a+ٞA��a��>�����˛���+4ބ�_�2Y�['�����9��=�n��b+p��='"TT�J4�=j�a�̐�v>����K�y:߾6&�Y6�ᮞ�i80; ���'$*y����B֙EB�P��B-;0����i���U���;PLB�)��3āh���J��������=p�9�.��͔��䳴�<�:��}|o����wd�s�Y�K6;��8pX>�v�[Nfq����`+-�<�P�1 �0U
kT�{p��|�XXHB�4��r#��ͭ�->�be˫&����;�G��M�k�
0x�5l�y6�x��iĠhy&	:�d�U`X���S0AB%�����a0-��R(]�)�\ñ�V.J9�Y��}};kE�6{	��p�k ��;��cn�%@��e�x�@���^���8ڄt(@�
t�����T�_��,�a��"��1�CI0���(De��Ci �����b)I_�����d�d	�<��c� #Pt��ls��!@b@�.�x��!�5��iJ��S�|C'����S��0a��k����l:�f�
V6�
\�uێ * y1��S�\"M٣�1���J�2�W?��8�	��4��@�Up�3}+��Q���JP��.����*iLB[Y{��J�q�SD���N,�t�{�Gу��� �����B�'m�`�̥2O!�ތ�}Y��q��G}��u͓�^љu:�ĕ��;_\��<�w$n���t�M^Ϯ8�2vE'���1VO}��c%������*{=#�넔�E�� ׃�w��qu>o�� �(�r�����!����ϐ��^7�b����ǾH*Ѳ82�B��DC؄>	CxN= �uj����=���~D��:9��e��yF�Z�<�b��|�%��		<��� �����P%wG�"��W����C�$>���ʟ�@[+ �#Z���1.����3�W!�|6���ctI���c�m��'��`�����Ga�l0G��xՄ�.�[�u����QA����Ba�L�t�N÷p�I�$8��R\X���|(��I;s`9]a� ��X��+�$Q9&G��^�*��8h��+χ� R�R�:Z��s�l�"�s��NSj�4��� , ��� ��<���R��������J$���M��� 49!��lر������H�5����pwS�23��GX�wH;�\�RI�!�8�\�k؞�c��2b�~T!�2ws� E)��B.S�CG1~�����r����	� �HE�����8u|�o�q�� ��D�"����_���=�	z"G�i�A�t�(/D)�r�˳9���u3��l��4��$ZZ�-�lC,0goI�=p� ����̔���2n�aq�� �����n�Z�g�r��d�|+S�Jz9�֥(<�Η�ǹp��
btp�`�6����8�P	k�j��"�<<og{�I���|�1����:����2��L���C� :�a ��b�R��|.�(�k�Й3�r�0Apg���rAP��V��O���� x�r�;?�/&0mzq�0�Q�7$��=z^�k�{l8�|���J4�T0<���IG�N��O�	�'��(!8�x�8*h:�j�h�2�4��;����C��_Y���Œ"v���Q��I�;���`��$ud �#tk���t<p�h�kޕ��Fz��tX�h�4�tZ�H�uE�
�@��B,�| �7�������q����KCZsM������*#�.R'3-��<wؤ��HqA�K��3�y�!�.��ʄ�K���9.�& ���p!��� s�3x�u����:nD鑞kJ���sA�0N������6���d'�AbpV���pO/����ә�#!+�}�|�n�P� `r���vW���˵��\vj�?z�8�lf���O7|2�Ck�xLvC/_ T=���� �V�!�(���@	<�s���',��!��>��8o2+����	H�t����ʅ�j�|`޺�,�B鵇�l�;��,s��o�pk���3?�|�|�_;�51�FLz_\�����l5��xz]!>���&��yB�#��uO�s��H���2��˾�80ـ|�������OO|���.�D�s-X�%�L_��G���77�E����׬q0r���Baa��λ��P iւd��N`S�U;-�����ج����|Z�~	�J9z�^2��#��BV�tC�au�Q���.�����>��0`�(A�{zT'�F��������.>;Lt�A�CDcIH�4�R Y<�4���u����6[30�3�i gE�y��\%IW� �'hm«5D6��D�P���Y��j�J�Kh�,���s��9!�5��r2�(2�I��H7�ľdN�a���ƾ�
T�X��aЊK����`XΩ9��g�8�J(��	�ܖ*�T���L�05�*Z��^��n��:��le
:ł�G��]��"�~<Y8��.c���'ͭ�54S{�}p#.!���H�q ra�eF]�l��?r��R=��$�;y[�0�I���G�!n���w��9��ǲNo1dyhZa�v\¤���1捿q�[�8�Bӡ�ӿ|уl':�����6v����ˍjv(;�9�q%��6a��~x�����O�\�b�V~�ƺ�bm�9�g��r )�0�gv$�H��,�"����w���(����\I��9�z�i�� j:��.B� �q�`�~AM;����*<(��x�Q��������d���W(���m_�8�Wc�� ���q�.�yk�&H�u�'�޻��T�۟z:���#\2޹;R�L�YE�/�1���V��0l6d?��`��� Yfu�2N��I�<r>E ��b�@�0X6"}�r���ۛ�q#��fL������Tv,�)Q2�!ǘ�O �^5�<����)�=�L�|�,5��&BA��	`+o>q�cB�v���/\��t��Qr�;�,� 1#���[G>#�X�����-���M�����%<;ؐ6���S'�#({G��	�X �RKӽЙ�o���)4xX���<s��	�J	��x�0>�P��6W�E1�O;1��IޮppQ���ڿ�@F$�^�R��hX��4�X����
�Ղ�+M��e'%D���Vf �����1����?�,褬�9�J\�a���|q��ۓ�����YC����;�F����z�̠:�ٝ��AIJ(U��!)����\��m�m��ʿ%*gSj'�y��O0E��b@G��(ab���ܺA���9���Ũ��+1��oJ|"�s��\W5��O�f�4d�i� ��UO&˽`�57����� ���� 6����H�zz�Hg�P �|&'R��#L(��[G�LC�0j�T0�����%������9��΋���\�cu]|q�Z���s�8l��`�%#?�-��:7QѲ�����ƣ~��R�/W�w��q	~A�|�hpRv[1�r 4oծܣ�+
����˼F�J����(L2�,?�`\H#>r����.�a6�뗥I?��犌�ׁ�i��U�Қ�
���\@5	7Md�_��Î��_���aV���y�e!#��/��>z����8�q.#�,��p����z`�8@��@�=��i�ِ��?\��d��=�H��h.L��5��E�Q+<ġ;˷H9o�
�u��&������3�y�~�?�M��z��.s� ��5uc�	��,9L3*�?��8�Հ �_Gа�띡�E:Bt;,�H8A�M���:�C���U`���0yE*b1��y�z����q�h3�u�sl�S�l�6�� 6�^�i�)+]����a���r?}�r� }}��)2-��1W9cp�l��tA>��VITP���+y���؈������,0�<�A}������ k�'� X��Bë��j���\gJ��|���UA��$�[��TA]��`��uŰ b���'A�w0
�j�M��LYS%��{ÚS0T)�1�M�;2/7K�� \����b��G k�p����Ѿ(��ƸU�>{�@Fϕ�?X�k=�����8ރ��棐�����둘��"���7z�ӝ�+�3ڹ��� ?bq3�s~�iu�bE�ٚɯL���ῴ���ő�GN�.�@m�*̀v�8#F:H+�x�+k=&��ߎ	���C��V�ɂ��@���3Ѷ����'���o&�I�
�ʅjt����C�/��㣡ۯ��/���Tz�d!����<w! c]�N��1��o�*8�v\/V���9@�)RS�G����8A�2j}�(f�֍�� �70 ��pmVR$P��,D�2��r��:9й{@ɝ	N����M��C�RܼO�� �	��.<}�d+�X,�b(�r��D/e�D~�a�3 ]K���<a�nT�W�#
��ΑH���Ҋm����gA�g�d� ؀� ��|{�]�ީ��#��y�~{�|��������� ���ŋz� xx��6�e�(D��+��k�PUH��2l��q�4�D��Cs���;���{��)��9���YFd���5m�A��KS�aELWr�W뉯IH)���z�2�����F_�5ˀBm`|a��#
��2�x�'
$��(��ۋ�Id���s]��3#��G���'b�{��V0�n�^�SF��N���a�AЮ���H�ga�:��z
������p������M]�������P��G_ę����/Ƕ��Z�ۿ��ձ�<YX-�޸8gu7��^%��E����f�誗ʉ��*��\L�J{M��3���њ@�=��p0�^5����8��s>R*��En�%90�S-�A/�f�$�1I��5煘wg��p%dT&a[ld�j�t>�]�p�� �X���&;��'�e��[lӌ�^��p��M�z��0Z�|�q����$-��X�E��u�s;o���寍��)J8ף���7Ň����<'A�1���N��@h���}��]� ��_���I�%�p������c׮"�����=��ʷK�e|qrC[�����y�]�WLV�ě�B� ����pln�{�� '��[�b��	��887���szF���@��n#�d���_[x���=�Kپf{����,��8&F�!K;�d]����.I�(��$hxޚ��� �8)���W��mt퐗��մ����щ̑�Zhm����s,_�I���Ɣ\4�Lx�F��l1�=y�r͖fc-#��[K�1"�T�k�8�=�̆;�7�5�^�˟|�r����g>=q�4�:�C�ߞ!X8|�����&)́�(�Z� ?\$�0�l�q�NWoT�nq�s��+4h���\xe���9��0zw��#apt�=>׮�7�x��8�����kb�"g��ҡ�J� n4�Te�YӃ�x���1�I�_������/���ѢW'x���ÿj���
��2ݷ���n�>r��O#�J�Bhg�8��@�SЇ@�Jd��5���b�l�=�($���k�,�<�����<I
��QA�5ŀ�,���=���y��O\�m�cICD�rYQ�Ixw��^��;mJ��iG���5S�Yr��k> �m)~%�Z��S���qj���u�Y���R�=y���A
�`e'p)W��J�Jd�STER���ű��n+�0�S"x�!�jlHL����<m��,G�2��r' ;�5���K�F$��,�U���&7ː8���8u�Nk,~9py��rz���5�J� �:;�� �*A�&�z�mm�5e���<ei[_(��۽����~�{��V��6��<̅_|V|��]�x���@��q���LV2\�c���o0DĂ�v}�p'�h	�x7Ώ6��h��x1Z���x��8��%[��yg� �q�� �4?&�Ӓ�R�3�G�l�{ذ�ɀ��o���W|L؅��KW��J���w���"��{f�^�d����ޯ_|1H��?�;�I�a��=���M
����.;��� _�F9���.Mb�m���Șf6�K�� ��R����^�+3O�� ����:s���"��M�"�:H#gBu�6(�ۊ�B��^���#naZ?�N$,��n7��<�&ItD�=����tJoT�OO��� T��z�u�Ɓ�c�Z?��&L�+;vu�OC�B)���_�R�O�qr?h!����̩S�h\¯�CI��� G3v��ի0��	�`��-�����N	k�g�xP󨛪y���u�po�.�*����h��\,�>C�9#h�=����c���Y�6d)q�ċk/��$��Ynf�|%)� O3�p��籠H�:�(�(H�Pf6$� �� ]���?�.���0��V�h�+ʄp�s"����&�%ie�\�\#�Íf�B��V��im�T�+l"͒~I�Vp�%g(�1S%��):>�cC~~��Iv�>��X����[��Vԏ��>����@3Å��ͳ_p��%�!� Ĩ��p}��V�7�	������o�rfo-p �㌚;/00�n��r���=���Q����`&�>��O��|�#�����i���� 1�0}����8k$��q�8�ϫ��C�q�)�m������^y'a�|(D�<�B��X��qv12��v���te��|�nd<���r�W�.J��o]1�qӼr���+��YK���@ r��y���$ِ�3ݎ�V X&�\{�s����̈��\|X��7��PD+|�\=39�²S9)��� \�2_�O����i@yX��7̺���\�8;䂨&L��?;��D���!|K3����X�,�?\ɵ����|p���	"�vj:��à�� 5)��A�h2��f*�	��Ze��r^�ʁ�V%��9%���ɍ�@�n�EoN�����Hn�X��д�gY�x>,)�ڤ�۸Zw�F %Dp�F$P���kL6�lM׆��/&�cf�/S�b@�<�Q/�ʂ	J��b�Z�^A�(��%(�Un�z�K�T���@��#�:�[o.@�2i�d�O	�V��c�j��|A?O��NL���w&a�䪯��j\C��c��-N���WL�M\f���ū�ǐ�1�c8Y���D(P�Q�](�%���k�-8�z��9k����Ǣc�ޠҙ����Eī����3Er9p;ut�:��ɢc�s!�>��n���B�6jR?\2�	+zf�5�"�
VVz��|�Hj
-�7B�'a]��,.�װ�ȵ�
yc���uZ>ID��>y��{Ɇ?����3�q4�
�Ȥ��� K�/�@E6N�lw�����!Ew.!��Ê<�M�2=x�u: ��g��f�k�"��%1$�a"\j[��ۤ d���g��m5aC�)���3u*&k��`A|sL���xA�*Y�A�=q�(�bt�G|�r���7�Bg�oho�5��PD�2�]6Q'��R���:0O�"Hw����"�]1eq��޸�
 V2���Rs�V�����Oı��5���|3'������oB�NU��t����nC�`;@�����h��o����f0�n�Gw��⾰�+��8�-��'䳋�kZ�T��x������A�mP{�3��P�U�2"�t��`\9l�+#���Ti�=�Y�5�2�!_]1�v�`w9iᯤ!��c�Z� ��z�[
x0A"pxT�� �R��D(Vw��6��"bP�%;3~�P
�ec0`��k'�Ě��kJ���p~{���p�]=Y&��A_ƦŐȠ��M�"�DP��`# �,"H�pPÃ�xF�Ø/��ƙRZTF
NU8�2vhQ��b�h2���Lo���IF�oj	�h��Zh)�`���)�y�㜫`h���,�=F�>��F�����g
O����6��_��s �G�_��!\� �!����N�xq����7,l��o3�I��f뎑�W,L��i���:�s�3����{_z��ٕ�/h���;�!|�l������������>��Hh�JA����{4��2#	��'��"&-�)��3��a���������ԏ��LfFnv��� jUb�xW,�ď�{*�B��-��� y�A0q����?�����O$p�G�$Yk]�Fx�J�����Jm�٘'���x����!����o��O���Ap�����Pه<b�L�R[�Y�c�.�Ӕ��� �
c�f]Ϟ{�vX�ˍP��\ؠG�ѓGd�)�.�|�`#�\�
T6&!b`\h�B�;nkMf̙w���X��Lb�M=���B oM�u ���P��	U�ĸ�/�\�af-�Yq�N�lv��p�kp�Z�T��,�`0#Zy(���y-u)"(� "�p^w�Z�0Ps9�}e�/q�� A�&��:�4�7��4��dm�D�24��]k�=�&϶�1 \ ް�J�����%�$L~Z0mذ�qnD�'�6 ����R���Uϐ�UC�arn[�*v t�t3���,�y�aۈ�L�)��I3�&�k>��s=���$�(�s߾b���˿�H!;ȓ�Z,��~8U9jԮ�{��
J���Y��'�v5�?�'��I���e~��:��c���ER�c����j}�c����0���9A�&�똑��Ӳb��QM��ٯ̜5[_�=,�CΎ���񩊏C��o�u���!(�R�@f8�!
�-`<$f���9SY���9�������W�s�>yd9XC2J\8�j���g�r}�q�� �N�K�y�a�ί鿎@)��ɾ�7�}��� ��pPK�'��P�B-����QI������xLI�{�h~E��Xni��9B�f�]�i���I�j��<�%2�ڵ?|�O����Ý�A�C ��P����5h�yLg ��S�����Hzx�8MDɑ�����<�T��r��Ώ)�6zQ��?��5� S0Ͼ�_<;0�S�G;�e�mp�&��`4��H� Ὡv�z�-FVl:3��A���D���z50��ᆅ���\��\�4g�Lg=y|\C;�,�Ν��B�һ���s$	R�JK�pHlg6���	5���8�2.�jP-Fu���e��"��!�"x����,s�Ď���5h /Ye� ��T�dP�0le��I�8��)��0V���Z���|b�^���:L�B�U��R�g��5�P��������ֽ�>�7ӧ�r��9�-z0T��3��eq�T)r�Y	�̥AV�2SgO�d�"y��~I��^���������� �S�����UA�Fv�m���	D��}}�S')����/%��'� �|]�<�����{������P7����s��z$�4�!QWj��AR
b�2f�9Z�Ŭ��� �N`�cO�l��n�la;�1s�v�|e_8v��vD�����#�WՊ��q��
#Ng��4�LO��	������+��ٟ֯.�3�,�,a��,�sSv���5c�8�m���'��6��:��<�ZD)F���3���w#�ˆU7���13X��@�i�-��޸C�S ��:�ʭS.n?~|p���'F@��Z�:R�0�xǞW�y3?"������~f����9��'G�=$��M�C��
�|�Xf��v�c^��Ì�!��sl��N�Jj�	U��,ۂ��,k �����LK�e@4ɔ|�U]6����
J`��0KX�d��fx��gB���@�(D��-{O������ct�dC>��� `����u���r��Q��
��(gM��HI��|$W�q�(0N Z����1�G9
i;����)ӟ.#�r�\À���L&<B�g.Y_�h*:�H�o���\���z� ��lw�"\��1ǃ��@&���<�Q�" k�\��Q�ZRL�����U�L�C4)��:�`@���:�?3B����ZP�@X5L���%avs�ӂ%$i�{��3�`|4X;�ZArp���hd�g8���Dh"h�Ə�[�j�P{�U3h�Q�f(b�lb�Kk���E�Y�U��V������ܟ�u����b�o��A~���/螠�v��h���d�M��J�s�C׋]~� �L�&�L!#�4�	�S�c�	t�����xy&V-"��;��������{�A�^Y/�4τa��rvI�$�ޡ��{?�u#�?:ζ�i��X�'����h�,����7tcB=�g���-�'(�W�A��`�AZ,5��m�E1�nN���8n�.�{�;�������>Yw���|?z1�WgZy��uQ
�#�RV�)=���_7RW��4�����.q�|˘� ���ahZ��{������a�yL�ȝ���-��� r�g��LV[S�ݹ/�����s��u�{)?����Y�ϐr�]�ZL���p?0��(�tF�hN\3���`p���M����u�/y*]������l]�+�'вc�?��/�x˫�ؗ5Ǿ��e�8K��	�xAOzP9\-<kwÑ%Nד�9��9;��C9�����U��ң43��M򂌶�� �UaO�k��}p�JG{�M���F����KV�/���|~�(n���nWN���b�T�{̰��	���c9Lny� ��G�nM��7 �ld� g4
�������Ԋ~=���(�6�ц�?[u���zw���2@Od�Q]ؿ���٭+Ǹܝؽ����^�BQ3, �t?���h�����w��g=��HS�>�{R�mڜ8�v�^�wc�3;�X�vB�eۮS��v�i~k��73Sq��̈́�Ǵ��N'�E�!��;��8>?=�t��`Y�k��!_d��v����	C��H�m�,����j�Ƀ�n����E� Z߆[`U^X�4�?�
8�Pl��"�[�Sx�Ώ���(FU�
=�&���1��r,�i�J8�=�؝�L7�4C�5�vXc�2m�,\	RlzkJ�x�4]m{�P��E۸gi�Q�@'e_�홽u�AE��x�/(*�3��S���7`_y�t}��s�ZC�5����!1�`0y�w>�6���຋��?��C�3�Ll�RL*ΕB��j�Ihҽ��y�~�x>�U3\�n71�T,��?���ڭ��8J1������܎� ��J��r��=D��b
�PܠB����Hҧ�X��?�+4�*����V�f��XQ�P��z8:������oV=n�������aS�n�_�m���R؏�=p�{�-���b��ܹz��'�����g�+uG�s:�T�������8�r`g��b�7�I��dHv��Q2��}~�2Ȩ���S2ڜ-�e����1���o��\���a{�T��s�et�礏)��a��q���g�|L����O��(pe�P������c�B�Η�
���ڬ�7�@�;�P�T�?�e!��7��d��~�6Z�.����1Cp�s�Cq�Ib��<�B6����M��T>�Aq��wx����ӟy�W��ɷ'���X�`6�PC�����S�(Q�!3�-�#^���u�PP ēD��/���bP~� ��AC�֭�Ԍ��_�V>�q���Ȟ�`�o@G� T   �;��a������ ��t6�庳�4�ze��I@� ��F$����^^P����4�P��6����tɌxji���8��;�/[w��E�I�>�/�i�UW��i�K��5�9 �+;dc(EkU�W�J�e�D~��O6��/��?�ݥ>u�{=]���EWh���^[��͊yAq�PYk�^�����Am������A�ڬ����bs�/����mXȹ[��ӑڱHz�4�p������G�~w���b�Wz-��{�E�[Î�Ġ���O��W����g~�7)-��+C��ax���Fo�y������·���e��.�}L�R��z��ѻ��f�t!��*}��?e���;��E����Rx1i���{��Q-�p{8>�U�X��ћC1�IZÔ����z�d��tA��e������gOv�)�w3��4�E��}z�G�Xy�f�'F���{׷ˏ2�0��\��F��j���53Bdu��3�n �U��������_�H�Y�_@����=E0����	��]{�e�Ȅ�\��v�� � �Z�l����W���~"� �sM	ߊ_M��?�؁��h��E�Zq��[�;X1=��l�k!'v �J��	Ă�[7�n�T]/�>uLo�.�A�>~��wT��:K 6;�|2�b�cP���u�����x'c(c���Z�_5��"�A�x}U"�ױZ��F�c��}�a1Gf��+eV����+`��~%�rn��N3Wk�&ѕ2��L�#+��~�<��V4�����$�[��M�IrDt�x����+�{q�`��H��2�#E~��^������;�Lfs=-��q�3��-�)��k]�RA����oL�.���_�͛���n�|l0����|�m�=�Z�Uҷ��یm�vs=��]3hI��w��C�_���Y�@$*�͙#�3�|�;}0�8&f��[j�{��9�&�=��ý�C�(���m荶4���|z)��,��>�� ��kr܍g�G�!�Uֈ!��!���g��$u,>�jf����/D�$�_�U�+y�q55Af�(�'͝��`u�m�2���� W��:h8�]���t�<6L��A����G�W�z�+���a�n���/M�nrvz���
���Z�8d&S�2�U��@`���s�1�E{��i��'�O����K���o�u/�ώk2V�v?����l#�اiĒ��L�����ݙ�sH���Z����pq?b�P����n���Z`���!<4�${o���$�UC�N��KQ��C;�7zDt;,��*n6�}{g�<.�X2O�=�����ȄY�����Y�� ��`7ǣЁ�?�y1k��8�Q����H_��٦k�� ܲ|�g�K��ɵI�7�Μ�R�&��elӨ��q�f���2��G�%�	�:v�+�+5�?�с}ǫ4� ��\��Z�)u4�l�OնB�� �?�s�E�g�OS$_DZI�d�`�a�/�R�K��	����|�sU}�'-q�t-0ۮx�ʆ$�L���=�۰�ύ�.f�*@��Q7�YaD#t�<�_��ʥ�և0��cq��QPuT���"q��9<��Zd�9��S�F7���4R�MI�����=jɇ�6�J7��z��j���=!�~��J,/i��S�	Tg>7%�¬�c��a�w껅aT�?�:��$��
P���7�X���JJP��}�\�{f�Χ�HΧ�2�%���v��VO�ug�]��;�
����CS����2}<�6r�q��l(޿��7\���Y2e��0����R!���
�0n�]��|��T��H���,#]0'��G�CS��o~4�z���q�"ny|1_�@�^&�Y��N�K�F\���72��� "��;H��Mu}�E%��Wg��K5o-q�����4��Wiw���f�>��:m�JD�����9-e����Y6O�9w<,n�	XM2��2>;�t�o#e�^���T5�sw�/�m6	/|����]���u��M���  RQ�   �+�jl��VT��m��	\���%R�w��A�[*L w��M��B��?���3���X^�$�b�R��c<���u� �sf�B=�
�F�=V/M�����6CI�������7����;+�α�д���gy� �n)#��>߿�J�0E�0�N����.�Vӄ����&��%Ϋ�E�):zr�R��K:b��z�u�$��x��Уxol�?���!3(G��d>��.�G���q�BQ|��NIχG��k�����59@����~O0Ö���������!W�s�yc1�<�[_iFȆ�r%�y<�V��@��v�l���*ɐ+$��_^�XlN�w#��%n�Hm��ɷs+
�[~!n?��?:����`�/>�߭-�����G_n�^[�OX��)x*d½S���c�!���S� �������g�m���p(i��u�v�����:�&F���h�.U�t�
5�����+l��������Ҳ�ڌ���L�D�օc=?2f�N�f�tS�W�B�.m>����ٕ@ۏ3�t�J5�8^^���}�����s�����V����>��+-������+#�t>Ѿ�Q7ڡ���ڐȼ��U#\�n�_�B���w�q���?~�>�}X�{��"��-�5]��Ffw�o��UP�k������,���y⣔�W�uu��|s�@ԓ�����੧c#���f�:��?��F:j�n�џ˷^�j�2����l�1�
(g�6W�:�`@��n�K����lu�<Զ/_����S8��8�m%=��v���e�7V��f�G׺ztk	 �q���vQ,"B�&;������m����f�D/��y���]_�(?�i���Q0���S(�G���!�UC��7
�3xY�m����	���
�|;bjdR��ec�����T<o��P�M��ⷋ�&�!���t��3���&Q�}�ʝ�a�4�9�׮�C�hؓJs�Ya�鹌�b�{�@Q��%`�ēcC��p[*)�HɌz��\ژ��*��?ݒ)�wU+�\����MחR��S!�Խ�h��:9�>_�_��RLH��s�j�f���^m@m��M?k��P2J��z|����D9�.��E�%lS"���=~�Yl���k�s���h�拭��x,�d#��M��a��+��y>4N�P��"܏��n�,m��Lvw=f���N|`���n���#@�H5Or�LS�8?���\nj��O������(kY�B��6%�>6!2�?���p�H�Z\!Nt_i�U\�:k�[�Y����e�l9��To�A�`YP9`Sɾ![$�?�|�d�d���qkN�'��;�;����{p�B%k�ې[9H]=�~�1JMC�|�9sFq�[�{�~���-�[��M�+�R VZ��ß:��Bi�p�~��x�@��UUśhZF9�g��$WZ�*�J$�3�
m +��P����>F`�тX���ի���2�4	]E�a�L��=e�f*��1��'䒄�YZ*��k^Z�Ƿ���rCln��h��EGNШ��T������4��?��`y\	JMY��f4�s���o���q�S%+��jL�#2ݴhX�r�`dk8�W'��L��Z�6����p:� j�s�����`��8��w,c���Ð�O�%3�=���y��n�~u(r-����oQ$0����h��ՆT��|� ��sb7Ц��γwAZku����7�>�Pع���d�~�d2*d��E0��"%��6�\L�ߋ=b?�*V`��B�b�Z7���t"=�t�~�%u��VK��z%d�C<�Xq��n Ru����z����O/��B����/F`&����!�M�/�ߦ����^G��[��wY���l��--ol3y��\��b�uW?�VC;��9����3�=oVQ��NMc��|xV��/�`����O�J��9@Msߴ�n����=X�^�3��E,�L>�?nQ,��=��_��|wJ&#e.��.ϥ��OB�V1�
��b�@��y���e�b��pzSɡ��5��=T���JK_���/�p|� �8�-/Z����^���?S�Q��o�tp�p�b��p_�4/�����WZ���Ub�v��� �E��'侜�ĳ��#}5i�r\Ntخ�a��KG�eotI�d��͑���r
0~���pB}�Ʋ@ɱ`N���٠���^�5�g:2���Po�<�A-���E<1�{<i�X~Z��9em��.c��He���SQ�Y�і�nXI���hP�yjK7���%�F���n��8Q���F�*����J�lnYw�b���)q���"��W������Q����p�L�x}�3kp�y�Ǖ�������5�z��S�-7b��e����M1R�j?�ɬmk͹�&�(��e�\�'�ȍ�\ZL�� �Ä*R̹l2L[�����:m
O�O=4���|c��7�h�w+J��(VqN� lѱQu�8�g9a���'K����l��m��L�yG���IbB�?�c��r��hϠ�j���P�e������7^����'���!Qv*�U����mA� ��v��ބ^<��& ��J�����#�ﺎ	���c��^C����+c��#DkBV���ѱ'� ^��)f��E��~O��"�c[W���iA�qG��G�Z����(�����a���ӹQK��_^�YU����;o����\c������nHp��a�����wJ"M���0��%~�f7l�2��X�?�-6�_Z��9�~�%��o���_�k�O�KCN���k�E�K:�,�|�7�˶G#LT[�S}�O��@!#G�ku�Ʊ�crO#���	>J_	��u�s��Lj�,�ԗa�H&}Q4�/t�Rھ2Z����ӭ�^��g%�`������T&GLT�G������'8����O����|�K�S�� {o��j��Fd\��/S���b�Zh��"}�XW~ 7�!Q����`����= 7���^�횔ρ"��~��/��b��Ї��������=�h��X7�~3�l��=�Z9wR�$��d$�ek�eBJF��(�U�^�2}�k^��Ql!�%���բ �|�v��Ƨ�n4n#�J`�!��Ȗ%��g�s��ة�!e�.��ue&��;��9�����M1�(lmC��AlG�8�?v'tҠ�Q�#���ɻ&�3L$�B���|�IcXw����	�~�擷����$��|K�2������kv9���ڣ�k]�:���!���C��L������9��xύ��JІ���)����%SqG�S5�z/��?��٭��(��j�kRC^!��ua;�O]]@���W��8�`��]M6�F���/̨���թ]���������{��:s	r����4؈�������eb�D���3ƒ���7:f�k��ǿ�^��~.�hQx�*��$�m�m��ݵ�8���r�I�F먍O��,��x��[�uH\�y\6�!���#��~\@a)<��K�T�3T�f��N�� Ͷcf"�ѡ��2$�����m1�	��5ߏ=[����?2��]
u�zE�� IRh�_r)_|b����ǣ*(���FRV�0�y�ᓀV)������K�]X�vB�E=H�9���4�$��4	�!�%D��5�s4�M#g���Ƃ��Ұ$K�]��O������Bbs����'
��J�oh�������*����O
,�J�?���%��n�ߔ7�R`{hLrA-��R��1�ά&��t
I�K����9��t,����r�Yߺ�C�򊨝��T�)^���?$���C�ϛM_�6 H����E�%@�*�����'���N�B����ٽ�e�l�vx���⭩Q��K`̈́+����#�Q�7���l�I?��[�J�扱��H�~��� @��KI�tUW��E#�%�بHu3>��AВ��o6qw\&�}��'|bc�={S�֟��5�C�0��뭈�{w5���½�)��|s���Q��K�9�I?{(��zغn���Õ�y��Qߟ�s���~��5^���c�BwW/�O�B����Z�]���_��Js'eLZ�7<C�Oͧ߂ދ�m���`�O�V�w��Aȧ���7f�sK��P���t���*9_i}Ѷ�8��d}U�ר!UR�`kˬ%I��r-�*J����?�3����0$_=>8�x���l�%/a�Y�$W]WK�[�g��_���#�[����=(�FYQ�xK覺r �hl|I�3��/ՄXmj�N�@�'��Wb���	�<Ƈ[��7F����&�ϻ�Xt������hȰ<Y)�F�
����\V�)�q��܍+��N�'ӥ�n>y�Ӳ�-�\�IW#f��2�ԉ1L���%��}U�hcp:E܀��Oͣ8�ێ�-z���LN�̾�d��R��Uͮ��-��g���Tp�3s���m�'�r������n�F�I�X��Ü�g1�úJ��A�Iä(HB{t� <���+7�ŶS��;��U�9i�DI��ݚ��ɤ��]�b҂~�/:`"�~�� ��}#�}��ĸ���Jz��l�50kI�"�g,����r�$�4��Hbp��j똕�5.o-��Q�N�NH';���1����[{��2j%���e�[i�0/��8��V���k%N����T�Rlv�s����gg�/U��J��ɑ����r�9,G�,e�"�>��
'%��Ԓ<wmbK�J������^�n��N��/���&�{��%8>�7e+�Fʹr-U����'����#C��D�m�?��|�.���5��F��~)o�E���P�6��F9<�uygI9����g5�v�Ds���.�_�*&o�.�D���C�de���q�������Z;7�m��ݖ�}g��+��K�M�k�����5����˽��-�:Y����ǖ[�QQ�ߔ����+�
��e�'�yh�Q��[�<zv�5u�4�?��ϝ�Y�H�����W�^���mDAm���.��{\6qZ���o�o�1���"��ѿ�������+�$��J��t��m�MT)2?����b��'3q��Z�۸�c��$5[]bmŃ(�K�D�RT�%����B�f^���r	�ZF��My!4 Fa�\�'�\8����O#���R��ҕ�Ї�7��������_�XBcG��g���Lq��E�۸��8��&�,�i��.a�l@�1���G�r�����GJ�����$�8�9>V|&���8L���
��p*��`�ʏn���!�Qa��NU�K�۲�^��,�ݚ��]�rI��=�%���jF���8�D���;���}O~N�>Ly:��9�%�V��ݡL`Ғ�����h��4ǝ+mo�
�S�?�b({ۏ��n�rY���v��y~�$][�@������4�ϛ���gl�~�[K#5A�|��_�S�_�s�=�����q�a�{\��е�O����7]�v�Z����	�N��U��Fd�4��V���t�U��io.���
�uv�}p�3i�{�J�;�.�#���J�CN��u�My� ��[�m�BX������u�oVX���AS%�{ű��6:tcP���e4�[:�����qӼ��h�R������;�/�ļ���rt���@(���v���k���Z<�e�Ϯ���~��y�Z5�Y��e�G�P���c� ����|:�b���*�����@��V	��"UBd�+�Y�2��hl�Q1=ʣ��w��=�)~e\d&��)lt7���.
$��Iz���&�Xo��uv�,� ���=4S$��m�9���0j.0{��8�Vd�����]�v�s�W9����B�u�!U��c�gH�e�2�U
�/�y&5��V����Σ��&T�i�����u�y�H��H�W{O��_]ù�v~����t�m��"SC���<�4I�U��::������n]&S�Q��0�ڍ��]���5�ύ��{]��̤z��f��O���:�Z2w�1���,$K�P9u�۞$��2�Y�9pO��/���spF�M��T��@������z���;T��Y㍓R�܌�4����@֨h���œ��X������7W&�ٰ_A��%J�J�jJXM��TrZ�|K9KQ��cv��[�\3���'x���%i,�:�Zv-˅���j�����WHyʸ�U��@���k)���ǌ�O���@4�a�*���G̎��}���x��(�V���H��^�w�	���B�1O?�=/��?��k9�ȗ�=��Hj�Kދ��ű�-��v:0�/�-��~ޯƛνs�[�Y�Of>������J�n��D?@YA_R9!�Ƚ��V�����b,���X�vHL^[���8��|-g1�x	�T����i��,[���*̬�B����C������}�^h}�C��YA��7&����hg���h~rB��'�'-��0�F���h��oF��"N�n?o4�aO.��8T6o=V�}s������g|���L��s���wvX�#O���iGK���0��B�N7uS��ܧ5j��U���������zGhP;�%�9΅��z7C�}��h�9y����,r���H+((*�>�yB����˞�+��I ��d8����F}1��1��"}�X&i���'�)�;�_ߓ!�2��yT�5+�Eܡ���������=#^Jl� ��C����P�v��)�T"W�n�@��&�仏��3���S�7��w�U���~��̒�m����8{�3(���T(���3��_�K�`����̗�dd_L�������<7\Dc#���q'+��Н���#��M��'�=��\saHV��0o����ܨ����	D���g7/Ŗ������׸P�i�Al��e_�h׋�mJ����0�*)W��Ӫmt%��s��Lp�K���/c	8Z-\�FT�&���bm�}\TLԽ�q�����7�2<@X�_���	���9�D�?&4���һ��ҁ�o�����n�.YJe
9w�=���S�����!vү���P\
z2B�^���|x���3(5L�Y��E�8pj���E�9�������ԏ����yn��=�¹-y��Q��̝��l*��<�j ��Wl�%T2(��%uA͚�f�������m��*��Z�[{�e�y�.J�\�#��{wy:F9d%o�9L���R�UC5 ��W7���Z�R�}�?��ɳ����7[��fU�4�������V%�HR�;2�����Z����ʓ'���0-�����}g
�EA��osu��G�y�7q��h�x�Ȅ	Z�@���,O?&���Ԉb-�6�������v�f�I���D���nR5XF�l�}��!L5�p �BZ���='ƶ�i�x-�nZ�#�8,b��:7�3'�X)f�e��j9}����@�h�5ZV��'�d�$u#h�1F�E �Q�_�o���8`ԑ����)�M|4|�*y͝�)|ں��'��rI�B ��P*��KN�,^ n2�����\��)|��>�01��r$�f���T�恒��.,bb�w��<ڱ�翈oeш��U��/��鰠�ܼ�4�j}p���l�(fzb��<o�����}����ww��]\o�#�Q`i����[F���}C_��*l�8G��X3�$^��F�҈�x�_�������+�o�W�l��Oj�|�{�"ɟ(����S)S���4�,�ܴorh����_p��Ɩ-�@����n�����O2ډ;�Iv4��A�D9��{��8�$��9����i��¤�� M�X�f2�}����L������C>����Q,� �w���f�w�J؎q$�'�;�@&���?�ZYI��6$���8*a$&y�A�-o��B'�S�pt��ނ�[>���4S��_]G�cB�:�Ԫ	%��m���~��g�^�".]Dv&�\��;k����M�O{=�~����	�\_PT�H�5EE�_vV�;��\s��
a챵p�)־$"0�;��3�T��j��2Ԥ��s�?�\�����]ϖ}(��t�Պb���r8����o�vM��+M�l'��n�� ���^~�!��&ċ�����ka�ͩ��9Ri$���6��`��!	�,���8�.�б[# K'�u���M\�b��%}��:+�N��~8(L�=T������/kL�6����ԏ��bp	��.�Ѿ3{ƮR�Gh�����^~����i�;��4�0tt�Kt��ݼ�0vwj�j=�
+��'�3���K��	�����~x`����4�T����qe�����Q�]E,�t0��Hi�Bk���Xk�
�ƻ��@�Q��Cճ&F8�ؒ@г�yց��NFtA=�	2�&>�K(�$�E�Dx�p���"B��ߡ�(��]���Ia;���dݙ����r�J�2I.�C�{�r��A{�$Ceț�4���\��P2$,$�W��EO�<�&�#tW�'��������Mn`��T�3��Ό�I�o���5mUG���&���eIaj�JZ��.#
������G��F(��p�Z=�n원��#/3;ϣ&mX�,����3���-k�S.N�l��0g��8 ��ׅ���BW7�g��S*�W5��Xz�'���D�����7�/�E��g!�hp�MN-d�M�N@݂���C`�I�yYU_U����{����Mq����e��T�(d�[-}BT����Q�~Tc�2���^�9n7x��ɸ�G�M����|wt��aX�H�*3s1����P|v�����#�}�P<
ɯ�i�����HG�1�z�nJ�ϏW_�N����1��x���=��;���A��0_�2P��cխ&�`� 4�e�Z=�-�栫���w�Q�س^�b�̛\$���}�: 3���t.�����p�-��"ё��QH�m�ͳ��ر������\JAB��]���MJ��	�1RP�ů��� A�֞߯"�Z�`�K��]p��P��t¨�9;�[��j;�.�C�����\�e��?+�����,O�R�'����%=gX���w���>���_))�3�����j����ם�"��A��!�{�0}�[1w����|}�Q��%�G�[��y��+�U��O|��l�{ ��tc@'E�}����3�U�gI\�cD6����tm1Z�\#YG����W�LR��|,�a^��EKJ��Y�9܋�Ӎ��2&i߃GF�����P�>�(X���GI�Y5Nu�w%R�#�Ϲ*aثk���;3��կ$�U���,���}9�N��84]�ǂ��*m����o<f�I����:(*iVt��R繱�1-�/������j�2`h&�\`m��2d(�>����J4��������:���� R���x&�����[�>Iυ�łK��[���j���Q呀�Yg��� ڮWA��xc�g�$����b��<��֠'�}�+�j�,Lb����f�?��Z����|Y�����j�Pt����J���(A��;�5e�R�f��2k���f).�*����Y�^\�s�Xۗ?4���5��ܥ�O�����Z���u��H�T7���RA-��yV�y@��P�tw]wp8�����T�	�F�A�w�"/��X�6���N�%e�=h��5b�*|��FF��W�o��⏪w�:=�+OC_|;�T�fg��=<	�~ׁnJ���[�W�yוa���FN0O)�zݚ�r�����Yp�1�3����� ��!��[���}j�"F#�� ڣ̈́P�R����ѥ0��H��?K���o��]T@���G� a>�=�����un����5����2�|p�t樾$��y샿�&Ё�1����h:�������֛���H�_O��!F8m1v�C�OB���ٱ��M�٭�͵�J�y�L�N�I�����q���/{A��=��v����SV�!�L�JB|Υn�|�9�>���x���h*?�M2)D���B��my�I�@)��zM!��n�[�3,vy��P��F����oyt�w���M��g�A�՚���J��"F��{�X�	�W��e��I�_��!�����P�V	�a�|��� )߂㏹�b"����O��35�a�O��x:�c֣ұ���r�R��ۮ!'o�qr����U��t����N��eb�[��S�.Yxq���b_��EP��<p|SC]����QcT�h�wDA����-�����I]p!��Mأ����6�5�\q�Cl^w�X�B".k]����I5ﵶR�[��ldҎv��Z]Vv,R��q'��wO��q��yW Ī@�/�B� ��S>��ߦ�<�[t!x��E,��R͔;VٟH��{�?0����@�9���3�%]�r�a��40fR�6�,�ն��Y	� L7������a��AZ(ar*3�c�P�@��I?Ė��ܢ�Q| ���1��|ӏ��`sml^2 EI:ٙ�k�Øf�ڀ:����yy��hӵg#��=�eTҝ�߉s��Z��T���_��xh����pmK��2ws;J�C��W[�sk��6���"��H
���`�t��m׆�8�aJJɕ�������&���_���$��1�u�_�.ߤ5<bB����cv�E!�z2V9����Or�D��31Pg�b���d�K�՛ٞ�k��t�E㤪�+�-��Yk>+@šjR�!���O��7`4 P�ʻ��)n�o��V�͏�wF|�f��3�7rEvu "wd��T�:�`�d��A��m�O��8�\&û�i%4���Jj��7���F�qל��{����u�f�0�^�߅y�.��ɯ����1���%�jps?��8��@oH��-]�����2%��gn� w4ny�O?���qB�9��k�T��)`۷�z���Q?����=Ωv?U���I��!v�ۦ�����^�~��4U��ͪ�C3�0t�Q���	;?/�o|��8oU��U�Ҍ�iڏ�%���L��D��Q�HƟ:�w��pC�زs��Н�1q����t1���Ljp��事|����P-KC��tQ�{.]��5"��d��B�ΫG�T�4���=$�u�0I����Yɓ�P�D�����tܬY��4�KEė(���$�;��iN�hL`�����&\��Nd7[-�q-qkc�i� GJ��X]5 5hAQ�g�d���^������m�(�������߯��0�v5�~��{�n-c����6����" z�Kë��&.��)_r�yY3�X�$!E 5-�L�U��i#J�h_�Nq�LGE�c����}�8#r��#��q8�w3�����?�;�c���~^J�����Y� ��OSR^ 3�'?�ywgC�c��s��/���&�5��g�5�t\F|P哑�P�Z�y�ã���P�t��
�>��rh�t>�a�Jh���8}Gt����
�Π^�c��7V��,���Kl㶂&��J��Z���:wʏ@��d��Qc1����`�֡�D�p�>��1���Tԏ'Ih�tƛ�<�v���/!@x�h����	v�k&� kã�Z"�[��b�m�Z�m�����:�}�E�]�ͷ�lG�TgC��� ���BP=��2{3�M��F������۷�2�W	�� xXt9�\�t���E�z$r#MK
�2'k��s�i���1C�z4�vE��	 ��Sl�l���N���t>z����]��z�[�S��{SG�����/!��q�qKX�Ium����(�_��U�A�F�޺e3^7��U@zR|u�6-e&2��EQ����H��0�fdr]���	��򊦵3���=d�GK�6�<���<�Q�gg�2K���5�?+EσtZ��/kۢ����#�I�j�,���[��!-Ԙ{v��_ZM\
�}�I�1�}�(*�#�b_ K� ����B������������rgH��k�\�I�_T1�R�xL�����۫��Б�����J���ă���� �d�Bw�Q�'ZKy�a���TD�	��B%Ŝyu/d�.˃���畨�k4�}z�&#��	�]���������<7E�}�3J�->)~Z�%�� b��+�l�gsp��X�������P�v���?Ƈ��)�XͣD����Y{��5�D��qх�1�^�7���>�F��Jݏd��c���>���8T��I�y���H0Ҏ�Z>1p2���蓽4`��Y���H8���]���{�C >��J�������>q�d����D֧�|�C�	i�!�$���<d��g=�����G&=�~���Q�2r��k�fB,
�{&X^j���}�5�(@�0$�S.�2m�P-�����(�#����.�",�Ic�6�q	��e���-�6K��z�|�-�\(k�N$�`V+4�!�rt~7�NS#GQ?X�>����zsbD����4��H"4`i�=��!�n�҈Qi�%r��#f�j �5�=]�������;g؊��D�����g�x ڀ�<@ÿ�YNIz7,Y�w8�ۧޤ�M�J����&"�h��y�$�-"�۞� �h��)��0$���M��詘V���1��Ҏ`̷g���&\����^����֥��8��סDr�G��^}*@���=oy�d�s3>q�V��Cy��:����ИU����HB�Z�]q�u(D6V�ɋ80x!3[~Z$�~K3���F׸���F#M����������&Rbo�D4{��P����w��k�zPb��5���R�f��Ql9��8E�+)�h?�N�.�^��k��Pd��j[�FD1khz�\R� �:��7���&*+/nԎ�߶T��G':�$	3 _�HlQb/�m���6�l_��}�I�jll䉔�Jc�o��]C��D<(T��9��(Xܲ�OOz`�Y{G]164ҁYĀ,���\Y@31͋e��uBG+�߬�� �XǈbsD(U�M�,��YB�E�7-~�K��@�G���p��=�ѐ�`����z%\sI^���i���
��� X����p�A|�������D!�E~<��]v��È�x��e����s�b�),���y9�+ �"&�=�""~����E��{�^)��.�Fżth"e����K%��q;	����J�@`�%8XfIt&Ë�8-JHL6�g���I%Bl�[��R �`�b%@p�/9���/e�E 2�$�6�к[ɰ��I;f���a�Xu�LLn�I�NeU_ж9̉��%�_-�n%���E�l�����<Yu>:Q�̀۴Q���f� $��7���{���8*�`�6���V0�&� v��{E%Xb\�Yݹ� �L�7� ,��&A�
J1��샛<t��%��1$o�vI��bI#}1����a��Ϛu��7�ۨ�>��O�0f#>jK�U����s�[��|O����\�d�"g7�����l���9�t	K��,Ki`�S%��M,�X,��e��1��Z�� �I!��9�zEA�'Pv�s@Ga��ڌF�[ףXA �3g7��"ꊳ���Oz!2�^,�� �NQ�XwP9	������Y-��ng�y�(�uh���pBdaB�$=.�7�ݥ!�	�NE�@eK�oN�n�`FaT�b�O8�ؐ�9�]�s0�$���s�IA�����L�*3"ɋ��-2�[-�������`��I$49�����`�Kc}_��X&�)qԾC@�9e%2��r&��a �A���u��� @����['�#�*�+ ɴ3�L��u�U��B(�RWmSs�sޒfUn⛵�2"Y�i�a!���� �|��ock��ш��r���և�!+"/�>K�jnE( �����jE""	l��h�L�VLO� ��&((/���Ԕ H�,0��)A��@��� �*�L����9���A&G�v2\�@!�B�L��D�L �Ф��>*x�̅&6\��م.�%$xpn���
0�e
�u��CE�F�VEr	V�Ņ.P	'�D��AM7� =nd�:�����S�n�6d8�d�6n���$�,��@�4�_wi?�I�޻�ZH��B��
t�m낖Kf�TܺDLG�(��"l���k�Ӂ�I`��D?jf$Ǵ���pǧ�^�x��,L\����&}3���ϹH����}�R2e�b�K�e0M��GL� ɗ�)��݄I�J��Fҽ/��1Q4�3�Y8έ���8wf� ���myL�^?N*,Jbs��4dp�Z�mo޴�����oǧ4�8P���׹�(Abrd��_� P��E�c����2t������%��d��O?�^30�Y�_�
���� 9���h3�K,d��0!j�S3g:�7�5n�4fy��` ��8 ��#���N#,Ÿ��j��u�w�[�h+��+�}TB ���B�n�s:뽜P���S���H>3wZӯc�9c8q!?�P�u.㦎�7�vh�L�o׃֠���&|t� �@����,D�l�
Hj&:���Q1���
U��zg���A��^�$�!o�� ��-K#}����DiA{��Ni�T����:�Au,^���H �/�/4Ś���6�١DKt>�1�DM�m����T�V�tk���?C��� ��&�ώ}&��"�ţv�����L�m�5��%�v��̑�ɥ��Lf*h��%Ct�.Hi[�]�rn�b�4��Q0H|ˎ�&P,�qg�!0���*���}w�ԡ��37�f� ]`#ؔ7��aT��[�;C<�d�`2���".mڠ6�r�"�ߵ
l�:2܂S[AzE� ��;s^A�+�}:Ǉ�J�%���;m��c^�5�����/�����grqS%3��C�S���Vْ�ŗ3ڬ��.� �Q
����ૡ'u6���5*�[�z]��Z5��n'5�8�q���� b�m!��X��E�JM�,G��(�-ؼLpt�`��+�����RT��7���ӕl��N|���!�_�ͭ@���bCQ{z�L"
��Ǝ�p��Y���LE˳hfD�Lݵ��m$m�C���b��;s�ߵK&C.4�����҉�;L^� Dl�@�}ҕ�u��%��L��lzb٦�I�T:εzP&P�u�-4N!�c�:��V���z��^�b���X��A��M�?�ʴ"����z��M�ƾ~� �۳')�xfs�����_I>h3�FM�n��㯏ߗ����{ۻN�WI� :�Ԡ6�����FEj9��Ūh1� bLn�&�z��>�%��ʜ�����D�� )ec6;=G���엎X�v�X�!��t���)$�N����[K�wb�3zϣFŋ�\���Q��;���n��\�����t�����I�D�O��I�-�������[�_���	@s���K�&��e'��ȗG�"R����s�F�{\�fԈ #=5���p��Ŝ���a3B�& 5�)�\�����נ9akm�M��2�����8�z�I襍���YY_�����<𴨇�~��Ԓ`û�,��F!P��š�Fqw@�%���ȋy��� +�bu�\��He���.��mg��6N���P�L�L_�^*�����H$�ZL��� �5{�H:�� x�J �bz���\�������-9�<��L.�V:[7�Y�Ի����j3�7m��P�d�!;�*F�����(���Ә�� J�F��;P :-i��{�,[�<Y� ��I9���L'o�Fh�2DO��|1P���jD1��=�A{z͑��7�[qS.����(�ۿ7�n�9Hǽ��׽+��Ë��	�b-m�y�����~9�L��3�s��R������(X�L������سc���@U�Ř�=7�U�Z��z�bF�:����TO�+��/J��&z���R�%���:�6���V����Q��B�I.�@����|Z� N g�ͦ=�\Qۿ���/zҜ����Xؘ둞��t�bw7�[v�^^�	0o�y���������%�kz`k��m~���1z@H/�y�+:� hm01ͣ�|U�Mg��C�!9n����(L��-��'V�Z=x�r�BM̫�w��}p��'�	g3�Jp�16Y�w�r��I����[��18�9?��C3 �ςƺ⎁��&ݞ��`d���0���Bm-�2Z~*��_ی��,��qoI� � "帴�7ǟrd�9�Z�7���$,�ɪ$�+���W3JRe����t��*�c�|b��oc���Mrm�����h����&�� �)F�a1�0²�� 3�Y���J2Jf����5/��Dɑ���Ҹ�b���֙xI͡x�cun���L�9�|�&bW��R�0��j1b؉;�%��������!f�1�55�'v}�H@����%B��38���L�F|��ỉfnn� �Ș����e��	 d�X�oӿQB%�Z��33��O�x�9j�*�s?����{��$���n&Y~��z&�Lrg�E�S�|NhB��� h�%ԕ�o�D"@�'��&����\&�z���N�[��^���+(	]O㧚)�	��l�� �s���=)�H���k;j/2��zQ�Pf|�����ݽL�eqA�=�����J�t7����6��j�[1��J�v$��"�{n�W��B�0����{����r�QJ0�9��X(9���m���a��'�=�p9����c���Gd��R�4`����z)�[9o���(��,��^-��o0z�9�
Q������f�s���ڋ �.oְ���}[T�N"~�ڡ�g\Ogޡ�^� �dy��ʈc������x��g��S�Z4y�B\��wJ�
g8��ϵ@$^oo��Ә���.����W-c��m�p����3�սiB?�I7(�{b��IM���$E�>�*	��|��[��HLR���[�4~Z�R,]�!�C׽��q�c��������I�-'��JK���c�<R�-y�KIB#�ݿ^�!��3�o>7SJ� ���z�g	=qI���5�89���ט��Jc2[�4vk���� ���I1��t������\�z���SXw6̬�-i����T��?���}Ш��Z�K�x�u��(l�����?T�VMM�Ұ䇭�^��o�ڒL�M�.��^���3�V���g�T�,����y��.�qg��ҁx�iQpcQ>��r/�|�7G|���HO*��<�� Į� b���!]�x-�x �]���q��\����uLz3�b����6�P��7���$�:�8ϴ���>)0`���8��Ă�z�Rо�-�E)�o������c�MZ�컬�f f>�;�'=�����a3����`asi�8��1��w�	��
z�l2	�y�fGC:��jar�����hl�}&syhs��b9Ǌe�=g�
����-���o.]�I��Eu����ۉn�V3�fzS	���3�+� J���zM�)����Ů�3-��N}���d���*��<��F���^��+�z�BM����JV�]j[	�=I�}�h����\�7���\�g7�g5Lw4��u}�F�v,���P��$}����ڙ��9��⊨�X��"^&a�N�Ie2� ��,R�{��e���ŻZ�]c!��Z2D�s�4@�E ��ߣ��}�>��/�Ppza�ar��;����K��⃱&�~�H0����ߥ��v��ػxߣBKR�{���H��v�y�ԏ�5 �-��m�Q�I��>������̊Amzb�4���~�-��8�L�E�z0�|Tۋ@NIY����Xr�� �)t�w�� �	��t�bN���M>�Mӈ��C������'�gz�&� Q����H�����j͗����D,�o�>���i������|�v{�/A-���=}?�30�?-!m'��S�R�'~i'��h��;����>>��.����5������	e��3n7>�R��kƌu���ޚ��G�����|sO{�s�����~�Ia�}��2��[�ѿ{�{Ґ,��c��� nv:Ң����6�5�����ݵH������'"S�g��|�IX� y�zo�>O�҄1%�<�`��q��Gg�A��<�&=��� �������Ü���L�S�7�6��3����)f ���	bY�ք�o�����o�7��V+}���V�q�����E�n֩�$w��Y[��>�-X�������䤫�����`��4�U�J� �h/���c������@o�����!��O�2G���ZlaP����N������4$��&�x��C��y�D�=�B.���sD�$]��I&�b�:�lwu��B���ON�L_�z���!�p���0�nP�e:�8��P�'7��f����jfo3�4���Q�p�x�[�F3ƾs4�L=��3$�f/�i z �ϥJ�%�k�6�[�s8��%�ןz����n���<Ǵ��R������<�w�g�M�w� j����8}�p���H�	4D�k�,R��Г����r`�ۯ�j���(��sw��ޝ���l� �wǂ����G��
�}��mZ�.#��#��nb�=9��x��ڜw�'�K%���1��j�g��U�z�����_��Y�6���,K���^�tD��>����PHX�)~�1I��|gq7�Z���C� �'$�n/���OH�8���b��u�/H��_�q�9����P�njNa�?]h��Y�c�hI�������G挠�X�+>ߢ�A� E>�T!G#�>�LÞ��萉�ܱ�g$��c�p�	������3��u���S&v�9��P#0<�1E3<w3D���������A�|5d=on4��HFv�ٶ�ҕd�rK~^w�T�����P�~u�޴9�GL�P%~jv��'�ې�G{��Ab��Ls5$N��~�w��3���FZ����=[D���5怜[lN9�%��ߩ@Yα;�\-���v��f��DмG��>��X���z�� H�v�v�W�K��qI����q� Zx���r�(2�߽4����T__���=����g����wY��6ϥH8fy�R8:��$�� 3DDI���%1��X�֢&$]?u�I1w?q�ޛ���w�Ea�Ɋl,�k�%�c���rQ��ө�pǜL���x��Y/��7�
�8R7|F��~a���lm*x���B�'G�s��Iܡ.YlG�Sj!H�K2Ƥ60�./�37�6�g>���Ky�CۼR�K��/-�Ҷz�>���f~G�)ID	�3�R��l&.�*"&�����I��c���ÿ��&\Zs��Hŗx�_��1Ld�uZ{��K!8-Ɉӽ�Э��o��1�ĳ�l� �,�vaB�9n��%�t/ޢ�y�✱9�O��`�Ns��n����4)&�ܙ���7f:C�*��ZJa�tI�F؏��iE�D���VI�����ot\�\��ח�R�]��sh��f0����w���#+>����Gk���.C='���t1`�[=��{K���x>�9��*���^�M����;����1HA<=��҃rI�hD/h���?�V���u��~j�,c<�w!Տ__3QU���Eͳ-������� h��N�|M��䘃�}~�Ytv��M�>\�0[���3REQ�N{���C�q��)b�E�q��JA��O�A	[�py���1Fed���?�����sgް�GVLw߽Ib�N�-��LS�\]Yi�	�U�s��An��G�N(���[t�T3+(;t��J�on_oh�%{���t�n���ة&�f��"�g���2=}m���Ǻ��ԗ�!Ԍ����( b�[g�>;���/���N�6����� 	�#���I��n���w7�L�cR�j����a�����d��.{~)���̛�+��w�b���7_��Ӕ��1�+����OJ�X�f-���^O�5�t����D-��� sZO_�� � ��f����x�8�\;��Q�=�.}3Qp��2�Q�"���BP��1G��L!{�^���?V��$�aʱ�hXφ~*]�{�=�Q���Jp�q#�+uŮ믽(l^"z�f�,��߬�Y����A,K���:���i��/��Z���~&f�=���XLo1� Lz�}�QXLDL7����{':��n��G����W���}� b�,��� �zn�3��&��	��S�6f�ݙ��$�ŗ>rV:A���_�M���ʊ�d�9flq�_�P.��$����[DD_	�h��u�	����ߧ��G
L�\��S�I�~��gP=<e���+�����E�Ú��^�|�b$�1ﾳ�BW1��x���*ɀ&3�C?�
F%��I
73�9�l�V�>'>��$,Ůǋu���KR�)8=f�b���m��5�����ך0 ǍK�iP,����Z������D3�0�Т��1���W��O4 )loW7�Q�2�7z�
I[v�hw♛���0'��c��/���Fi��(���>�yA��b��{}�Ф,+h���SD�;�����O^��� �$Y����@2�~qH`78�u�}Y8���e|P��y������f-�ވ]�������,�}�*
��H2O�sR:�7����g1�b$I���=ib@M�5�D,�~嚉��-���iۼ��\v�Q��7���B�v�|~h@��P�f�[��i��2>����!��߾N�!�oy�4�RǇ=s�֙�d���4c0�g|��'*yl���C�����w�<{�LM3?/�J  ��u�ّ�7��uC��1��n��"�h���T�9�j��q����o9C��*1)�d���₤�ʯ���(dr�u�@_��m�)%��L��� �%�e�/Abo�-jr�e?�HI|�-B}�8�V�,��<�X������,��Q�whKX��?U������FS�=oqE98̙��YΉ;Jl��i�ә� �S��^���P���U�[T��zY�gX���\�|���E��4BDǎ���i	�n�'CQKو��=(,	�o��t�U��ɒ!�����(~�ӈ�*'S�iL_�b<ۭ&�x8�^��-f��7�>�{���%�$�jo3b��o��!�ǥ��)&&g��$Ze��<�k��3��Q����Q�<R@�J�19� �>~���:�<b����i�k����o��� 1j ���朶�`@,�bO3zT�h�������Ď1l�椻*}E���oclb�� Q�M�N����G9���)��^���o�h������Ŧjې��g�ujheT1��n�D�L	������p<�=7L�(9뇵�U���}I��"�и
��î�2Q%oee5��i�N0ߎ�46	v��ڡ�r`?~�#�ء��gR2_7�R �ŋ���	{��c��*��=�F�R"�Gz��6���JA&2O�� � ߙ������Q�N�)�-�$1BM��t��r�D���>�%Pci}�6
Bm����R&t/w��	s�\�3#�� �h�Q��z�;�m��P���������FH�6�úH�^&x⮁̰�����a7�b(�r����eՈX�>��,��w��#9��3634��	���Ԅ���;��8��c��Xd���S��~�P��O���J(Izg�ߒ�r.r[/JX�������8q�=�B%������2�^~s4
!}K����̹m6�-�h���⬉�f#}�҈������K���`���ܼ�B���:��ޤ�5�����z��MIo�[�}b�\q��A"�Y���6U��bNR�LT��&`����R����Z #,��s� �'��zP4�"Y���K�(�	Ly��14,`�b/�c���q�^�$=�Ol~���w��1�J��� ��Y�K��1�0���(����l�PX�Y�X��X��Bň�w��	)"q��d�O�� ���� ���A�Ư������_u�����?Y�K�@���C��o���ͫ�n�ZD3�����.��h�=O������:��1#3���E�1܈�4�E��vi���q2�P��=kw�O��cu07�	�;�gu��bz��BXϮ��B�p���)�G��� g�9������F$�����~�}+Q��8�� 	�mϭ�@��fbE(g��R�<J�g>/H0x�)����cҲz��K+��*&���>�s��� ,��,��R���b�B�4�����jD��(�u�|z�
Q����Z�l���B��;��R��\gu"�~��G\t��X�ܡ�ű�Yf�&r��;|�` -�5��MC)#;�OX�v����^m�>��PI��Y�y�,@[GB�y���Ay���!)Yˋ��褩u7�f��5�������2�'&o�;40c��R��6��X�J	����)G33+���"}_u<�R�����R�q��RJF�&�z�( %�qlT�n�����ŉ�?������l�&b�#�}*J�	�|sP�/{���.V[ֈ;�>Y�2i�w�S�Z�S|߽�)`�3���eW����VT �N�ć�2b	���ٚ�B�F.�߭JE��l牢��[I��B������f�9�i�T��ׯ_ZC GӧCؗAŝa��D |ߒ��U�"}����)%��-�:j� W���wY&�1dˇ6���0Y/^y�r1})�tC��F�i[1�O_�i/w�g��D���ne���'��s�ۛSd��θ��qvmB���ҐX�Kb3�J�HH.�C�V������$�rb{�'/���`��6Cv��k�tz���vX����J��R��� ',�b�F��zy&<��9綽�J��.����S�PKD0��}a���`�8��阅	Y�� �x7�}�n֭�=�4��˷���ht�oЕ�aw���c=�x���LD�[�Apz��֌���敄G~��H/�� �{~'�n3�j9g�{z�9&q|���ir7':q����~�B&G'�59Ak��c#�3�
�ҿU1}�{��+��̷�NmI�I�sҠ�3巯n�c�ڈ�&��Њƣޅ��}���e�w�J1���'ߞ�H0�Ǐ��bzķq�n�no�֠�5�E{M�2���"��2�M�(B��?�\�7�'�Ғ!6�gYu�Q��Gy���l~�Lб3x�/���K�����p3đt���ϜsK8ɡh'շiq��*c��})֜��8��� �DI���*�f����f���V��a��8�Uz��� �P�d��Z�²��!bb�?�C ɓ(�u��=�Q�ZB�t�;t��%��y�x��/j]9��w����D;&?�0��z��P�A��7�jaR v�����X���৙��R�m�X��5���1n3�?�ԗKs�Ǝ��-����S3ߦ��ĝI7��zY�v�z�.����<x��.z��CDC8��%e#��T�����}�ݖ�:�FDGS��y�/7�b'ޘ ] �_}�e�qz��E��5�@"��|�S"V�Ƽ�^�8���� jCh_��K��%+�2�g��� ����k�AY�_>{o$Y�7��H,ק=��L���գ%�o��"�oؼ~&�bE'�X��3�9�w�@��)V�g�3A&��Lz��h�̥�;����l�zE$�^�_׭"�Ε�=�F�=Rb\G�5D��zE''9g�_ڭK�3'�(��L���BD�l�x��$lL��4�	�#v��K0؈�bb=�xb:sY?j�9v��x���|M�5�G�3hEn����ji$˒�:��L��$�^p_�Nh���os^W�S�-���g���IBPC&Q_ٷJ��i��-�֤-��� �W�0#��� ��M���1��343�r{������:�-��H�@��'�FK���Dms.��ڀ�˨�� �boW��^�g�i�#S��mL�	k�)�#���RR1��$��O�RQf�<qBTz|d�xZKnu��f�oބVy�37��Y�G{� �+Lǭ���L�ނ�-�M﶑w�� 1=k0�������ot}�y,u�"�����lbm���%��ܜw����3n����Pe���f��\Gz$�o�]�(2G��y�R�b9{Oj��C�1�+G�/�Z���~9����F�*�։��xw��� jH��QOO�*�ɐ;_T,��[_7B���g=;�% ml?y�M�{s��U�]�O9������ׄ��|Z��}ezI/0�U�|o���<��V���;��$sX(Eķ?�����a�ͧ��d	���|^�R��[M�D��{��LL�]�n���$�12n��K��I���E�����M�g�n�K�/��z�U����h���� 5@������N>Z!f��1�J�2��=sN*�I11������<X��݂��L�Υ���&y.g��\� �u�����:�'<�֚V�	#/`��{��ք��y��B,oN���8B=Z$��3���(��U����B�Q�	�3J� bm���D�n�㊲㫭�A�Lͧ�O��0;��ۯh��$�?�C����|T�S�H�8���ɂ2l��7<�ۏ�H�=�Z�_4e�	t���X��/b���o.c��9J����?�s~�I���H,��V�[8�Q�O@�3cX;��r�e�����S���� y���?|��A3=�ˉb��� �ȓ����^���,O��8�;��e��|_�N @wβu����� �)���Z�A� ���jw#��>jrݎmxqGbS���@Bo,Kx����@����E���\�3y��c�t].��آ������w�޾�ǧ�$V&2����=y/J�p�w��)ǟ;�r��CJ�c[֊"���E� [���Qa��K�Lv�1�>p�3�A�������~h ��1>}�S0��L��ѯ�������j��|Tؗ�c8�K�19q�҇:،?�(�?;J����D)��4=f3늒E�9��E۽��փ(,�� +�x��H��O�-=��x�J�n���"�ۗҢ��31�����U�o���C��'� ���*V���j�2��D�ږT��F�D^G��	�Fm{�(%3x������q��j�
�m�^~�����%t����uۏ� �e����}�3�^}-5"�����_�1d�>?�&ǧ���):=�ϊ�-����z��vs�x��?xᨠ�ǤTD��uo��T���}e�Iy��u��s�<5�P�v���=fh�F����&ݨ_(��_���h{C^�����GI'X��*A�z3#td�:F��qBI���-��d� [���\W(A^���5agی����L54���\��j��7���D)��R&َ��#%�D��-{\�4`I���D�$��8�h$B^��_���]��tQ�s?�# bك�\�^b�1kGZvF�q{&���y�.a�ޚIb$�_2U�nvw晅�L@� �^�g�E�S�w�]�&k��<��D���,Z���1�"[x�>�*F��s����>�����,��'�ǭ@ U���ls��ߛF}*9;�=�j8�Y��`��K	��Jbu5�|�W[a�A2��ߧ� �)��)�t�o���ͣ��nKϯ^8O���3ߗ��Z�>����)���g�1D���?g�a��۽i�X�����^��+�u3ۚZ�;o��#�f�$���������w�j��jO��e��#:��eۛK�|}R4z���\�x*�q�9�|50"5{�|߽�1�������TGq� i5�oxM���gx�6��/ϴv��� �l����5���9 ��^�Qmt�SD,"�f-��`��c�zFx�A�B6���f}^�Z�O�hI+���/Nz�S0�^�3Չ�7��^[�J328�3�F'���<q�ɝ�̞棽ƭ��҈�8�>��*N=u�#[���������|�J�x8���3@3�F�53Ϣa�� ��w�R!3jL�c]�ba[�5c�6��1N�����g?T#K�� ,�c��ͳ�����#��K�NnC��߱FW[��CC.b.��V�[��x���N	�������[�z��6�jx���S����^�0��gݤA��3��!�Z>��� ơ�.~��ώ\}�ǳ���js6g��X ���_5���/�]��|�o���6v��(Y̇���� �����H��0�1��F�_n��(�9[?�Ҭ͍܌E���O}f�;Z����@���1�׏֩Ӝy�E ��&&�`d��J�Pb��:pZ&�d������ߚ�p�z[|MB\���Yc9��@�7c�_�1mA���2Ù����ړa' x��"���K���[�'(���օ����ރiDOO�!%������ ڒ%P�0��z����Q�2����P#�F)Sa�*��7�z�E������0^!��E%����R�L��O��)ř|/���CRs��%"nԫ�NFأR˜�� *Ll�y��5i��ϽE��Y�� h��v�N(HDHF[��(H�{�?��&���F�l�[ϫH��3׊���g\��fZ41��{	HC�x����#���JD�s≢��Q��h9��8� ��/�۵8A"�1�Q�y�;U�t�=���ϯ_z��z��o�2\�h�V��`�Y<�x|RJ'	��ߤ��8�b�&���������C����Ϯ&��:G|O�$�����׏��P���3�X�H�i��jܫp�׉�H��.����Km��W�D��� ;T�s�XϥMbA���y��u࿷|��3���eu�m��Vo=g��طkQv�Je{��vc��E�.��$Q9�?TI�y��L�bwc��O7�I!C f-,�њ�bF�/yf\Ck1(�i����j@o��e;���IL���u �Cbt�n��V7�2��l�q�)�8!�3��J�(��ä��H�I�f{Ÿ��'�#o�s��΄�����Ѝ�:~9�B���(e�V3򁉋w��Uat�O�ޙ���h��2#�����2#"l�n��a�o��f��3h-��ҨN����/3���a��-ޘ���tZi�[��:S�x��Bc�X�V�x��0K�~m1�5��^=�
θ��#I�/~�P̓���]��buA�m��z�u�⭈��bc���c�^�hs���٢@q2o����P����&��a���P�zA~���)�h�y�Q���TL�Xh��]���ץ��C���h�l�#�v�7ݧ׽D�3&=��4���y�@!˪�w�l�m��>�ԡ}�� ��C	�ǋy�0���o�֔�+�i!iϊDoBL3h���_G��#՘�H1�S��fg�_�)����ތ�&�b&����۬�D�,�[�y�w��%Sg>"�����]&s��/&�_�A�3�,~ifbqx��8E�Ǵ���r�x�	A$�Z[ktbn�#�z��S�X�\EV�Qn� ��7��ޱ@:y������l����Ee�B�z���Zc�~�b��8��,@=;��-&$�Nq� if�)�D^?|[T����?�A-?^�PBL�if#x��� �ݶ֭����jb�_(���9�T&�q>��B�9��ㆋbݭ�C2�3��
�f���3ˎu�TH�O�>�����K{t�(�AV�t
bjY��g�H����q���Q���0}PPg��zP]ɜ�� žDd-��ie랽9�Hv�Z|�"��}�.e��i��ao��Jn�����P a�Ҋ�-����*݋�;����#���@.��.c}x��b0	`��5��֛e����B���\M]ʽ�Q6b2�q�l��l|������ ɫ��w�D�<
ϧ��HY!�D�e�'��h�x�>�N=��K_�lLE�@���[�~�Ej{�����A��ӿ����5|�u��I)�G�6�Q<D~���l!�?5heY{��o�5���ZTCn�3�}� �I�מ<[�J�A�X�T�3��=h�x�J�>z�-����(\����/���I��P������暍ff�f���̭�i�k�.b�RFh1�o�z����P�m��i�8����~��؇=�>� TвI�03N@e�f7��͞�o���9�y��	�wҔ#���A���@Q��?�$����(�y�9��)�9�~;y�O��H��g]���:�}�rq<��~jQ>��U�����\��S�AI`��7�U��c�Ԉ6���/Ϊ��b*DpO�w=7J��@�=���ٻ>��r$�&/��~�z�Ӿ�	]�<RF��u��O�.9")y�b������-�2D�b3�ޓ�x��B!7����N������mП�� ���K�s?�J%$���:��B�6���>��@�q�^oR �E��;�X�?��@�+�9��ڀ1���y�٩�;�<M��}�k�F�e�Ϭ��6�Ϫ�Y��9����~��Q��Z��3Q":c�	���6����W)�x�Ii뻿���R�L�?�Q�L���I2��LB#=\s5��t?T�E�f���v`�o/�z���:Z�����^��a""����o�{ޘ8Y�a���!T�����J3n� �S"��o7x�V˜OJ����|�i��(�g�.y��S��g�����?��S"Xק�Q3=s��;��g�pW�����FW����Q�9c�S	�����~�>&�l���*A��οb��=�7��J\�۳ҝm�[���7�w7-󚅐>��=b�D$�����ޖ1xz���ւa聘���RO[ro����'nsP�N�?�-�c�g8��YY}q��#�����g]_�n����Lu��j֞�|����� +@��>�� )C�`�"c��o$���뚛@�rk��<0�e�bޔ�p�ހ�@oh���	��ϥ���(K���9�� X@���q�N�i�L~�� )���(@����#|���6�e��BǇ�S�>)Xw��M�~�r	1����'�ՂC�`mSs���j��鳷�2s��O6�Wֵ~�jL�0q;���.s����Ҥ����r12?q���b���� i�b�\މaӫ����=� �v>�T]I�aN�P�Lo���r��i�t���@>�k9��>���٫�O��k�=� �d�x�S���O�~�`,�s��%�y��_����Zq>3�'� ���x��oRaֿx�0�+|�j� ^�"�x�>&��d-�/�@g=����w;sW*�I�3�(�x�}cژ%��<�.��"/��i�ނ��[9��,�
c<� ~j��8�k��V����(�<�hBӌ2��y�0b=�ڐU�;���7w��D����A�w�,-���#�i�[��2�$���~�����AA��X_断��_�w|�V���V���1�	{	��k
�7[7#�[�4@3 ����%ɋ7���/V�� Fsn���X2۞ǿ�D��q7�W�`ҿ�.	i�\<� ںАs��ǭLU��m���R�8����Nߊf�!��sL���w���i��J�y/�9��4�)y��8��/Hy��n�8��em���(��o5����6��,DoW�꜒#JI�}3�,����k ���m
a�xơ����w��H$#���2T����R3Y ��b�Xt"1����%Ԝ7e����z���z�2��u<�^ԓ�y��s�/�����ŧ�h�� �y�Y7��� Z��u���D�8ٹ�5o��3-I^���%�&8�9��9x[>_�RX�Ԣr�*���ӧ�Z��n?�B����ҙI>�ZZ&gX��P��ͯ��@fl��>s~:Q�Q�R��ʛ\I.�]�����^��3@Q�%��y�52TW�9#ҋ���c�����#�v̴sy�����A�=�'�u�'Ώ�EA<������ctXd=f>��6�&K��ޒ݆�,L����κw�f��"@����$���X���w1���1$���� 'u<º�~�:3,G��Vm�s��}Ԩ��~��� �F!|��Fz�6u�zJb{��⌦^��_�%���� o�B�}fh��������@'=Lyώ)e#מa�#�S���%>����Xm<��|��Cbן��� "8��G�Jz|�YݩB!��:�Z2��u>b&��l���7�����$Y��ַ�g����P����5��7�^&��p7�Ш]Q8q��/"u��ij3�������-�ni��%��Aj���� �:��1@������0�n[��]#���{D�1����q�4�z'S�?�9��d�X&�1���i�o�?4� ��&��7�Z�E�K�Zl��|7� �9�n�ןz-�\3l����H|�b���D�D��5E�Y�7J��~��C�}m�����{n�	�'�=���_����|P�s�� ��E�+x�����?�{���� �{��~(0NP�|M�ߚQ�'�V��~i7nXg�E� �us Dc��i��LZ-՚�Gg�����/�v��w|9�d-�t�P��i�� |�㯎�����I���B�.q�uPnUE���ZT	1�?��`굷�Зqu���QXE�$kw�4L���ȶ�Bů}_-JYd�t溕��5�i�9���Z8�:Җm�xo�*�g��~��H��gX�*���n��e�޾��8�"/-͹c��v��x�	g��7���bt�o㩌R�:g���kj<q�|ct!|~�>�-fY��m� �)��Y8~x�Zf>��(&������HL�'�W�C;-ex�b�H��	��z��)1�Ǥt��TD,�>��߭C���N:�,�s�qnjGR�����)E��q�A�ɻ��1V[����v��VZX"�w�ր�o���㭕�Dˌ����D��K��3mě҆�d.59�h�\����K��[�����=פlS�o���Z��ណq�A���G����Ƌy�ޙ����h%,�X��^��n|{SJ�\F_?}��%T�^'�I׮���nN�*M�LΊ�Yy��9������ �>Q>&*�,цL�s�� ʒf:{����҄�������
+���ſ��t�?{b*{Nyq�m�49nM>��;E(=�����~:U�<y�h������t��y����� ȹ�{��������g_; n�^�(Y���ËR8�����xֹ�A������$30�6y��&5˚���� 4S8?�n� ��f�#�(	�rC���%��*;�9q3oJd�,΋Np���A��|ɪ�83M��t�'���G{k!�o<x��gs3{}{P��%�{4F����Tdrӏ٤�ן�X��zv�K�9�EI����W�=xoZ�ވA{�u�߭#�w+2=�K��|R�#3�� Sޒ7-�d����R '�����n!�C����6��#��"x�*�|�'͢�� 9L��_[7�R��s�y'\y��Dt�,�d����L�����11���P�w��i# RB�k��	�PbM�ǌs�%H�p>�j�Yb�g3�r�Ţ 3����]��U�q���e��X�z����lD���(�!d sq9E��h�ϛ����yP��|�|{�ƍ��v��� ����ߝGZQ�	��3h��S�� Z��S.�/�H���<��!�K��|O����7%�դs�;H��JIL�qb����y#�ԫ:��f��s�T���fbc�ЛgR���!	8v<����<�&手a�o���	��{ԡK$�zpG���ج
/��� <�(=�ޕ��g֬��.�R�wY�؊��D+hӌ=}hLU����Jn�i��-��8�T@"��|�F�$�w��  	��e��Η����[T�ng�<�[�0� 8�v��W<���1/9���C�=hN�u>�b�}�tƀ2�l��3'�9��Ͻ66���7�#	��ϵE@�|q1��G���(R%�#�� �F�2��G\��2��N�u-�{P`8��֜1#�=3���,`[�o�Hª�:t�����ݸ���D�|&1֢-$p���v	9�!�3�c8������ ��ip�D���-� h��3Ǌ$���3�x��zL�,���A�u�-��� j�1Ƥ��4�"���	38Ȋ�$Y�,s3���S �dG<p��R��Kuē��r��h���շ�t�B ���&�b٨��1Ҭ ���X�
-Ğ�9�����&z��f}9�PU�f��|GZ(_��i��[��#ۜ�-��2�Q�o](��@��5���cקz�o��%�6>'�#�l}O��@`_!�i�H��|��RHI�I����P���������ޘ�k������{�8	ON8���f3؊�q�}�cD�sނL�1�@Yon������}�<���� |Q�1�-{U�f�t���#�3���6�u���K]��T!"9���#.��z�������)v��Ry���1>s=	��p�7��wR	{�nb<�ͩG��Z���M[���M�/�����<nm��Ԇ�M /���=朡����h�s6�i��Gw���	�o��Y����-��^�}�nϵ)m��*|�� ��,�.H��=E��`I͋��Yo%hI6%���你K�|~��3P�ā�s���T^P�I�<o����Y�r����u��Е�Z����z$d��-�� "cWm�Ij�#�|���<ԃs��Z�kD�l|{Rd��8��*#^[�6�x�
��q��L��A�� ]hL���c��JE�����$����Z~c�E�w/u�	C�G;���U������c�!$f$��O=i��:����y�`�凰c��	��y�֔]���t�����g+oJ �'�E[M��9��#N�?��e��_mA��PLD�$�y��=��v�7�/�o���Wg_oE"����2�ļx=��f�[a�@DM�/�b�����o_9hA�1��L��~�� <�5 �b'�M����y�y��M�-���w�HYK��if�@Q���~�Ñ����Z�E�E�R�-��
@��[f��ۡ���g�f�5P��[�
k�U�hTx���ٙ/�����X=c�|�,Hb�gY��u���嵮��
W	G�g�t��6���?���4
eqyq��&q�#��u��ՉX_%����߉�]o���P�(�8���K��G�׭QH-v� �>#ml�rqzsRX�}<������ng��F�s���~�X���s��O���sH����j��?��ތ	���Tq�"���8���⠳s��k5j@#>�ߐ�]<�����}T�ü��J.�x�1���M�z��G6�Vl�� �ݏkP��c�j��O��8�������ʐ�zGߊr��#��JH���؋sԥl8����N�ހ�[�x��p���}�� �ȡ��m��H1���ߥ2�+���;��o��������"w�x�Q�Sx��%�3���_�@���� 2��{�jdYK��戇���_��P�ܿ?�LУ:s��oߥ�RK/	����$��[*31�5bj!m��y� Nbќ�wH	OAn� Teh�����z����^�/����7J��$wX�p�ǡ��Am����������Im3�� �P�t��S`�.����女#Jd�_���(bX��� �|[����x5_�B���bM��z �C�G����c��	e�����)��^��g�QbА6�@���tl
��۳��w��U�df,�y��L��<u��2@b�O�S��'�I\�Z�6�z)}��[:� ������yީJE�1l�|ɚԾi�q�ٜc8��9���E�y�g�����M�5B͓����Ł�sk�|R��ō�ɞ*Y������7g1Ūr���}i��	�3�zU�~�D ɶbowTn�gNw������3M��v�z��e�O� "-���K:��߭4�SS��oN��Z��wNb�Id��������G�g��K/,/�a�	���HWւL��~ic��h��N^���X翊@����_��$�{�/4I�F�>zM#-~͏�e�r�7��s�BC��l���@l��B�Жc��d��}1���B]$͒T�f�Yt�Ǉ�Q�qf�P �er�v��o}�!��1N���ͩf��"l��3%o�Ϙ�6#!�-���_\�L��|�hLl���� i�!Y�_���	u�H�~��^�s�g�Q!���d1��4����,���>��O��M��9�����>�Qbt.����$���]1У*%gK76'���,M�wCy����Kl��)��s<����0�ZKH_}b���{-�z�%��'����D��\q�N�=�x�Ko� ��LJ�5s��BC�ӚL�<�2M	C�9��{*N'�	�r�:�hzTRb#�RL��� �"���R�i��7��ф���� ���0:���h3��TH/XC����1B����٢��o���������.�o���b$⬣��������%�-�k��r�o�j�Dru��  �=��Кe��}�+��ܥ@��q�=iN�gв:����(��'����!��6s�w�ac����b�6�%�<���B�ns��5��s�U1�u=��Y�zG�-��f�ffو�)����x�g��P4�07���Sc%f7=H���+�?bs�H"�g�?��
 �a��P<D�-�-���j��?&�犕$������	.�PI0γ�K�P��w�`�W2�f�|�L���.��b��ZJ��T�.���ũ���s��P\ı/��z��4/,����\�o��M�A̫f1==(%&��6�[���Y�Z[oϊ`�a����n�a��>%��;�J �N�8�L͞�hI%�5aqD��1~?yf���y��q�i�z���+	�H�ڤ3�J�b/2����//��H�b9�W���v��$#���(�gj��L�>���C �zQwƬ���t���@���⃔F2\�Eɒ�W�`"d���|�(���A+�r���T���ŧ]����"|�ܞ!��[&8$;C�ְ�\o�?%�����aM�:�|ޑ�w:ix����z�ꄒ���f3�z�2�=jE3���7��ޛDۉ�8�>��P�A����ޣ*�s��K0�^'8��Q/~��'T�z#i�f��v��?��"rO1n������w��Y.hg:�-x�EC@ٴޓ9�|"A��op���	(��=�5Z!���^���Q*ř�� �fff%��R�L���8�hB��}�Ϗ�W&�_N:ڠ@�
��~�P��D7�o#�l���hd��j9��ۅB˙�w�,xۊy�<�13ӂ��fq��:�ރ,1w}N�c�2M����ަqU�-b�G�m�K۪�q�8��6�E�PgZ�x�iX7q��{M*r�ėα��j!��烧o٣��)��V~���z�Ku���8�SY,�bd� z�ϣ�Օ�C�}�pb#���(����J��^��`]l��O^���q6��� ���ON?f��/촁H�o�u4���� #� �����h���o���-�Q�v�1�oL[�g}�zS]/�>�H�I�� ����W����������ӚY��K�|�$�v��6��շ�sS���8��?Z�R!3j����Z�>c�3�D�]�������)��v�c�h��C���|��gꥬ'S~g�X���J^ |s�G�Dy��D�����Ƨ� D�� ���f�O����Ce����2P ţN\b�l�=� eikLZ|z��Q��:�j+{b��9��		�c�Z�p��X�ӂ9�t}7��g�@�ˢK�ˮs��=��Ve�����K.%�w�����J�Z޾����<� *aix��J�q�αM�b7�'ǚ�${�^���)a�t_��`�8:��
�T�ﺔZ�O�5�&�e�u��$�>����)�WN?M5"'�|���V�'�� FE���ͨă���Y�f�������8XLb�����Ǫo���j��J�a�R$M�1�qH�2��";n�
g��ތ�4 ���8�Үq��b�jr�W���PD���QȆ&`���"%������l�)!���ak�<V��X�-H)HN�_���"�V}3ΪVT����#Yͽb������ƨ	�?�ߥ`�����ꢱcdܱ֠1�w���)��Ş��\B�8u� [D�7�i����"#>���%�fz���8��D"u��� ��%�2c����M�_��c��n#�o��	�b׋���K��0�p���(�#F�t���ݷKa-b\ÿ�B���HY3��Hcyr��g��By�]�<Y�!�L�<p��5fS$8���\��.����S�#6�f���LCӚgz�y��x7e� M�H! ��{U�ͳ���h��3=�6^#�t��� �-Ι��[ v/��N.)7���)L�o����	�c]��kf���8�?�B��/��P�E�>�����`��v�b:t������O4 5���y5֔&g�*���/L�\�}�M�)Ps鹎mK�.q�=����zU�D��<�F��xϵ)'�~VzEL00�7����� ��	ߩ���,��_x�����٧.�ǵ�]�u1������ λ��zd('�~hQ�Ź����F8��~/4f7��5r����R�{�ۏ���� Q֐��)&y��<��~�����@	��jH9x�Xgҡc�ٷ�UĆf��_t#i��;sVyy����Q���4��)$îY�Y�*ȴ��7�Vf���7��e�?u�DL5����"�s����2K1|�s�3A=,��G�4��m阾x���≓d���������S>P�{�2�H����ʊQ1������ݙ�j�����"�v��9��J=���<^�l@�s&��kx������Z"����b�)bN�-dLD��?������a�͌Z[�sA"a8� 8���&�?1N��3�9���Mg��4ab� 4��[E���2"cI9h�Dql��I�y����)c�7�u�.~��P_�=i�S��~��Ay�\�1�f��t��
ͻ� ��̅����Fͤ���� 7��|ՠ�}���i3��Qa�9]�� �V�q	���>I��^br����� )VT�cӵF G!�Y�^�m��?�)#ۯ�uiv�G��0���������^&��q�(�P�`��B���VM�8.-���.��M����4�>~Jd�{-��"�@�8�<�o��,.�����E͑%�z�ˋEﾞ��,ΖKNq�)V��m�=<�0-yM��x�YS��}E��6�&�/�/��
�;��❌������X��� '�Q�-)32gxݣ��HPX��ޔ�p^�����5���vC��XfE�����
�}h(u���[��� �L��6�������&f���K1�7<y��H�<>!jJ,xS�����ns>�ޡ.}cڔV"<}R��q�ǹ����ʯFO�6�#���!}�"�K���	b�X|Aך$k�� 7�@�}`�×1���@vM�g�l�K��w������4�NS���jIZ�`��x��]���&����U�="��Y���A��Ϸ�ô��[��y��]ə�V����=+@��L�T\����J�R#���Gy��ꞛ�K� �|Z{������Q�H�����K������I[��T�����W���߽K�����բ7F3�~�� �>o<e�bԶ��މ&,�ӊ���?,�E���1Ng����7��P�'���/�"����)��j�N�#=�S8�3�v�*�Fx��jt�����|]#��T�;��� G&�L�H�`�"c���<��{�(���.
f~g=)�V�w�o�J���_�gz�F�w$O[_�y�	LsṔ�f�le���P  Z&-�߉�_#sf�8<կ"l���@�������4!D7C���C3���H�&�	D��ȑK0ɲ���D���lf�h�7ue�R �d`�8l�-�D�3�_��$���{a�G0����-�p��Q�L�^Ә����T>��`7�Ğ9�bf��*y�̟�U�-�fu���0�����b���G��ūA�"��H�3�_��w�n�1�qۉ�"g�?�]#,E����A	/|�ϭ@L·�c��i/6yy�F[�j�ة�	�F;-�sS&%���bh�\�3��֒e�T����<����z�\H��>|V�#���߾k���6��h�e'N*o:L����ŪncS>/��pv��+ �/����pY��g�7�4 3�y�o�A�Cٗ�J�>Ϯ=h�6{|y��n�g� `��� �t��c3B㧌ǚ �������j&�v��d �����ﳵ�MHĶe�O_��@ Ʊkۇ�Z� M�I�{�>�-*�c2�Ɯ��囪p&�Ȁ�B����"��{N7l�G	K�':� *L�Mɻ8F �{PY)F�coǿ%��3�#�*@2+%�L-�m
ܓ� �6I�����o�@��m��S��/t;n�ƾm�b�,Bˡ[�g��e�*Gw��ɳ+��<��{J�/r~�@�L&�ǡt��ӱ��e�_8JCd���w��-p��>��p!n���@'�!�3>���7�lڦ$��m{Sǘ��ڲn�mH��v8�J�׭�Ҧ��{Ғ�ǧ^i!�S�я�|�\o�+"2���?��_'3|��$�1�����F���Ps���^�G�~q�S+����>*)���]#���#�3-�� ;�Tۼ�s�`����ݪ����o�@Cy��z`F"o��ڣ:Ý^j���3ѵZ�f.}O��h�>b��\�c\�|�g
9�_���I0璎���nB�2�k��P,��b�}iI���:��9<x�F��?T��� ��9#��ON��x��Z�Fm�:�h�Ȑ�$um��AH��K�q�ے���F|��N�uf�i���J���:;����&IA,v��19��� "ĭ�ꏓ��ZL��▚ԄY��n&=�i$� ������H�����j��4�p���w�����]�.@�l�C\n�|Q/�D�,���q4b�C����
$0��$���ʒ��$dۅ����G�ne.F�g�Qaz�Y��LG^�X�-��n����.EZ��/��� ��y#�T5pz�q�2I58�D�M1v���bژG<t� ��]����L�<^�9��˪@�?[�Ff�k}T�&�K(�ט~9����,9��f�|<��sD�[v��f=ڰa/G���%�""M�I2���~(U�=�]韚$^-�o������m=:�����7��}t��q0���s�h��m����yq��<U�O�Y8׋PFD�`�X�x�I3�Ÿ��+�h=ڄt�fi 	����s�/��\j7ۆ�kf?�!�#�|T	�w�mи|;���T��}'��>�V)��-�JB��~�j�;��zsB6Y6���� �(�}v擤��8��Ǫ8BM�� -�bB�#!���k�\��?���-��+����wN�go�|E!���,N1Sa���HGN��s���"���^�;�X���o~��*tl��N	� h�,3��4L4��\�NarI�O�w� �Qw�~�*���zD�y��1 ������3A{��)���?�R���翵"����k�) 'PM��Nq�f!�$bG��DA�n�'O�[eF�"z�f֗�R�2Ĩ��{t՞1K���ZK��������M����3�ޕp���� Ҿ����V��D�>��M�s�\y�SNFm�{�T&=����v�/��i
�~�֯x��0�䳂uӥ�(�����Ȕ�DL�7?�T���5�qI���� �`[>�I��5$�s׷f�'�����f�!O3η��&e��4��g��`�͹�E�u�l[��RH�7g��-��6���[��VRM���=e���U�^�� {f��eylg�[�"7�;Db� ��IF�<�4�m�!��3�0c��	��ͪܙ��2T�L��/$s$u9� �b:�k����_��/�w���/��� ON� e=w�6-�/~+ �K2�k�Z�h�  ��2���z)ĒQD��[�E�AC*���bՂ�=xr�-����"���l����@9S�6���Ү��?��B}<�� ���r+h��n�%�ɓ���_��}� ��8��i�(J1�s���-��o�b'�H���9!\��5N$�f�pg����������d�1O"��l$E�Ј�$D��'�"������4Y s�o�4�p���F:T9�M�z���CĻ��$����V�1��c��Y�%g�t� �ͯ��w�PH'm��*�,�5o7�,���O6��[��b

a8���c+h�=sQt��9���ߍ��L�A2�R}�g\���8?u;a�o�����G&���iNd��Tm�H�9���T�{��RF�c6��SD�I��Zb� �҆�����eV��� fb�d����ŵI9}ř�>h�[o��E5��J��?Z� �lrt��%.��I�@߽��D@e2X�Zԃ�{�QI��z�� jb̡��:u�B�D̼�����.��n�P8+��n_�]@q9�Ŀ�A��S��ץ�HƆf� ���:�Ζ�*�fs9������Nh��-=X�5�5w^�FY����N��_g��yH')������B���o�ֿZ�W��x��� C��1BD�)cN}zj�C"������"eDD͋�MsKsOX��W~� .�_����s/e�óQs�8����io��"6%ɴٔ�$b��10�/;n��&0i ��#?��i�Q'6M��8f/ˀz_���0"�㷭
�²�#F�3�&kb�r9�i�t+m_�-13��=�߹I�~5�y��I����8�N�鬥��Ԍ�{ʐi�'{G�JO���v�2ӷ�1�b �z��J��k>i����Q�y͚�1�>�-�G��ԇ����2�E�LO<����m�������DM Ih�s1�t�������1.4Ư��u��Z!�&׼�צ�t�v�G�z8���Q�g��-�Pk�C+�b|]ҟ 1d��ڴ��؝<q�F츷���j1+����m{��RAw��߯�������m���P��(	A3�zF��̾��"�1�sO}o���<&<���H�_��%.�<��H�kz<M2C�����'��5��Y��T���mբz��nfhE��怓���-�ǵ9X3�}p��6�!	�,���	�	��s6#x31�uQ������	>陱:�ľZ 03&g��a�10�p9��4@���1����'22�XV��)��G�����>+���(=�*s�hXD�[��E��}
o�Hgʒ��z��Gҥ�=������T���(��faZ�Ӑ��[Q%�Y��%���2��.��?�u�پ�ͩy������]���������e�w#�ҙ�Ī��]��FD:xj�����Po�r�_�B�HGG�S4���T* 2z����A|�-���*����!~z2p�D��4�5��NP�"��_JNH}�jt��r�{

X齝�n!i�:N*U	7�X�5*\����_4H�E�O����hX3�� Ν�B���?�rz	dD̈\�g�#�m�f1��d������,���� (��&�1��P"�X���En@��g5(z����@,L	�=�bP��p���b�fvF�;~��bx��AכߴR&#t�;���Vzfrf=~(n��Ƿz�����_�J�������=� ��3���xd�4uǸ&et�C7������l��d#��7� ��u�oI�H��㿟�
-,y/��B�X�1���R�$j�`\��;4MK��zM�ϣ� <�!?��5-��n�k���k<�mK�R9�ſ��dA)R�����f���h�\AeĦ�i p����z�gm�[;���� ���=
��O-�S�33u�� �L	f�W�A){��S
��P�0sg�OzE�w�e����N�x� ��� )     !1AQaq��������� 0P�� ?dR/�k���"+Z���:� �������a[L̲f>5��1w_:Rrw�m�����s����H��κ�Bŷω����6s˷�	�;_��z�>lI��h ,K6�K43����w�j`$_�ԯ/����آ��K����$��Ym�BA� lm���-��� ��Z�d��Ŵ���զ}�O��	I��#�m�i���ݾ�X���C��_��˟RbY���BLE��t�?'�/�f��6�r�+y�u�\�a���Cg\S�-�{���\AI��%D�� �K[�+�d�2[�x��]M��N��\�=E:f4��niE<�� TڐCp{�����랍C",0���(�W'�-��<&�%��Ɠ�R ����� g�)"�$�-y��ͩb�tF�Y�(+F�gdm�P��b�=W�&2��Kt��5�NIݞ�[����������#���K��GI�֧��3�J���i?����IH!��9Қim�L�عD�w���߮jQ�|BK���\�e��#`��R�7y�ht�혷�Z"�e3�W���^�rM��ޙ�ճ@o���wzf�d�gk��F�������g<?MCf�u�yQ����~�Jg�Apy�lt������mhU��TM�v�M������W�i-�M�8�o�����P���Y�a�{��n�EꠎY��1Ȉ\ؽ�n&-�:���$Ia��f`�x(J�ƫw��P,̷ݴ��&i��d�t��a�f��u]1��b hQqbm|d��0�����`���$�R�P��̱$E70Q�)2�l�;RH��L�Z�T3pHcT���-�hH�x��M����6�_��J7�gA��jM����\qJB�0���;�1IX�b�<Q�d�mhE�_[S�.�8T��%f�%�?��I��݃��S!�v�yر�N�	/v	�;J��{6�'���5��u"h�v����uw��Y�M�t"%)�m���mh�,�"݋2� ��eh��Ĳf�Jl����w��A1������͜��ym��qZ�9&��^�M���1d���/j�-��9�����"&w'�N�5���O��ҡW��Ƴ�� (f��H�g�*�T��r8w�k�h�ᾳ�*	�ˡn�����S:�r4"M�����y���������h�b-+-%1 -�
�Xڙ��Q0�GL�V�nP��Ɠݚr�����
L"1�~��!'Begc7����'�Zv�(�8��xސ�+t�e�3�:��gߗ:�쁙����3(}|��Le�.���y�E��A�zT
��[K��F	���b/�K!"��LI��4�l☡�L��?9�F���~zg��(A.�n��Q
"�Ó/r��	r�'M�2�3(	r#7�L�b*%�[*��H쐭�}sQ����t�6��i�0�\_�Y�1#��g]�4���ǮA�ތ�L��$��4XK���@K�9I�:m�t�r��}�K�^���v("B�W,�i��4�f���y[�!%��!�lR�!f��E�VBri,0�b�%>��bfX���� �P
��pP�X�����e,)B���RH
�ͧ���S�BL^ѥ+&8��M!��F)��'�3{s�����o! �	�Y��(��e���F���I{�$t��2�Ь�����kLv�P&$�s%�c��4���1|� �Y�,6p䃃O�DpSݐ��1��P2�Nƺ��`�@�2K�t��gs,*��Ӫ�W� hm�-���$d���jM˿^��5�C��I��'j^�k'��x�Jz`f���}�5h�ذM��T�C3,����-%������$�Ke��	��&(�+�$��bd8͞��`�cOI�2'b-|���ɚ�.��㊲�a��9�i> ���y�-�w֘����s��*M��� 3�ڕB|E6�@G���f��ـ0�<��KI��t�h�M@A7��^�e�ۥ�i��W������N(H���Ǩ�����_{Z;T�*w}5�Ӊ��g��OF���+����3,�z�5~�\3;�O�5̷ɐ�,Z3gKd���㯽P����3l]��}�b��/3>��Ԑ7��:{P��9�x�k��c.tD��Oy��"�et���;EJ��rcNkP����iֆ3���C�S���v����-�u"�a�',M���i�>h�����ҊP3:fOXN�^A&,�z����0�g�:�:T����Ys��6�;�&_\Շ�MW�4�mxXL�q�hP�$���W���!�,s0��������.d��]<4Ϝ��M'/Y�O�Eه��N��R��! c�,ϥ8�Ce%�����Z�&�%��
Gq�CrØ�oj�\efpŋ��� Y͢_�z�PV�i�9-R�	��wcJ�������H#75Hq�3J@�?hZF'��^�*�yjD���`���;o�Oz����Žj!#a��|٥�������d�T����I��r}�Ni������2Ria��٠E�sH��~1Jr�.?�3v�cAp�c1��I�Sj��G^�Z���$�;�H`�y���l�
�]���*��Sq�/���4�W�ey��@M2�m:�Y�S�k��o�}b���*��ٌ���2L(�wΠ�4�l0$��nv�@.��L��biW�8�~���A��I�Й��~��Hz�b�b�!;4��Zc��v�3�Kd\ ��G��!s�[u�؝1���%��9�������]��@��ك_�\��;C����w�9D��}ڮ0Kb}z��V�{��PfC�6ψ�-�&HR\oΗ�]$��6Ky�� �^D�zL�s%��i�s4ۉ��mΎ\7�y�dc0hk}})�d�bd��A#",�q�z�K}e�{~h��їa��Ɲ
p��cXRor(�.E��gVCf��@l�es��IA2rB��D�kP�-������Q�!g6�D2���Z�@�&-xpg��S�Խ��F5�0H�h�3z�0�\��$oڈ<�x&�8��P[3	�p�\A���1������`�����
��3�눴s�^%���W�N�r�ׯ�Q�t��L�-tpN-i���6����o�jM�\������.�.>��<��Dm~~���U�m����_ص�2"+�k6=3B@�K�O:��	 %1;o��\m��=(�:~�I�+��"�.uw�*d��F&���ɻ��i�C�~�h�6� ۮ�8L@߸_�x�i�Mٵ�<�u�yǢ��8�,�
8��H/� g��,B"_��G�E�u��@���xާj$��|&P��j)#k����]v��a��~�@$q��Ǯ4��H����[
 @�wv�@ܷ��bĸ���PD4#��>�hO"-���/E��|����|e��\u��%����z��$]{�lM�9�r+
F���b��[.��\q�T��%�6l�=�Ү�N���q�<���vi�ԣ$�b準y����t�{�O$9��?8�L[�Dm��R{�j�H�T�h�Ɂ�f<�a]� :^�)���$ƞU��5wţn��k����4�^K�tԘ��w�0X%l-6���:��);{LZ5�`$D�h�N�vM[�N�<P��6M�xL3��xf��D[T�۝��s�dr71�S
Q�fm��zF���wnfױw88\Άs���S����8�m%�X�ٷ��"ЙW�юf��`�>6P���"�X��4 :��9i'� �{G{iJ��G��$h�-8��c��RdD�{���ym7O4�(Jc�9`�n1�M8���&n ����w��$�z�M�M�Z�/7����:�x��CM����7q�aY��5#P4�N�y�%l�/;[zyP.pJX��F�����j��̆jK�D��>��WS^.^�\3m	��*N��"1�^볬k�c�@u���X�2�o���Q�� ��*@&�������52�]�L�m1pXĀmh�zx��&��o[������{N� Z�as���#����$$K�c�oE
�DB-K~g7 ,X�l�w�1�#���%�0߷%	:	'��u��j( �h6��H����3���z!&�1Lv�Xh%�ݐ��E�I9�� lh�b����8͊-�H���h[b��و4�b�
�$�"b�ZjL$.tm��"E�ld��4�:U���͹Ѿ��@$�.m�g+7���)3)\I{�2�Ր�X�����ݓ3>U�-��Q"NTJ"�獨̋Z���ng�Z���X�<Fm;�Z$�jeS��B��[�\��%I3|�f� �ȰC�k(h8���mh��f��hdo�X)aG`�y�F9�HBd5uC{1�M�7� j����8�c�����l�|��"���N��v�rFH��8�-�KG,�3	���������0���km5 T%Խ����h訴�	c��AŶ�[|g��4�!�{�։�e7�f�qpJ�.�P+7*UYv�ܩ���%q��_	*ɠ6���X�.0o��@�k3�v�)��m���T�[OޑD4�}qo�b�%v���ƭ��ƕ�����ʒ���Dm����@��1��n��d�F���ث�:�����8���]��۫���tG��s��l?W�#1v%,�]W�BhfI���&�%�C�j�ΛI�fiY �@a��-�lT�-�R�=�W����6;U��ai"�j����7�U�B-��dB�D�-�լ��#T��{�5�[ʹ�՘®M��#�Yܖ�� L�m[��LQ6�nZw��7�e�Hc����!KQPIa��Ą䄰Zw�j0Yh�"^�C�Cq�����������8���Zi! R�˞M��.9��9����D,C�}�Lo��hY9H!��L����L���#��*ȑ(,��5�s�bL3Fe����3`�{���{T� Ap�>[zZ��!!b���mSu�y�6�ޔ	�,������U�D�PۛN�T�L;�`~m+��VY��� |�bH�Q-{�k�@N�݇��PRH0����r�qN� ���}�i$\9��^g�@_���֩u	���bMC��&�����r��l�.`��Ck���xւ"�Z���OL^��������{�m	1��h�^rd��8�/Dk�u� )aS�\X|m5���Nx�J6��?�j@���[ZgH���\`����fC ��-o_�Y��
�%�}^(�L��y��љ�m���5�{��t�j;>�t��^#fw�1����3źS:�ay#1��ޗ$M�u'���R��q�Z��Q��R�#H6'l;��*�������I��f:[��U9�&��-�LH�A k-o8�"-8�?�oI �aD�,[~�0I�1�lsK%ֶ�ش�M$�����LD�WV��\��%�pG\O�R%�$^� �"�e�9� {�j[��-���<yt�[�)k��7�H���d���֝nwe��w0�ŧ3H�p��;ޒ�@e���Η�b"ʀ/�0���7X1c��#S@�2),��Kh,@��F�ݽ�UI��k�ѵ2W�0�l��B��X��S��F$�8,��XR'M���6Re�������NV��֝�D��fړ���
!����oQ�
��ʾR?�c!��e���L�R��N��9Ͽ���bf�9Blo58�����妬/6�䐼���j~Rj��g�n[Jw���,&��^�Z�X��2�G͝d�$yD����ބ�aq{��Kn'4�9��{���օ8#i�wҬ���3��zJH�O�ޕ��3�$�1�����Y>����%q�G��.�;q�ىƬ� �D=�������Z��Y����3'n5�c��϶N���ȏG�z��pgZ�޹��.Ȳ�1�sڡE4��� �o��qQ����1�C}K�Lg��R$.���j��ztGjG!�zǍ��C3�&/������۞�0��g��)Āƺ���}*lE�܋�E�j��anϒ��1O$��a3���.U��/��Fˉ��[:�mDE�"W�N��"0:f���-�h(݈�[�^j؆RCx�b�ϥ1�D��<ǌQ̉�K���.�H���>�d�EnX?g�M�z�^�QB�t	���n�1Cr���^lE��x�4U�2=f�HK�0t￡@i���vƈ��,��v�#�J��3gXݱЩ�z�hL}��U��,�u���	�����C���.�n2mκ�&�'k&f���|�����oMe��(��x׋�W[H����j#iw[��a7��bZY�6�kLK�J���˼YD�5�q(���7]/��dY�	 c���Z��y��߯tޚ
� X!-}�-��˖���68��OU؞�M*{r����h-��}o�jH��	�����[	.@�tj` �TE���-,Ep�e���͜F���~*@R��ȶ��2��HI6����b�a6��h��E��06Θ(�JJX�ͧI��6P��/ź�G���P�ۥ_�.�M^/�(o���"u�XL:�PV]��-'$zt� �a�}�0۰���<�[m~oJ�e���֘����\ä�췋ϧb(���2��ڤ��m�o�{���,��3L�H���Ls�5%���h�byӭ#,F���K�'�p�;�i�ý?9&C|k�MO		!ű`�Hu�	d��v��$��0ffH��&7��O#!�8f=�Pp�F�����& �	���}i�"`D���y����vF��v����%�-������[\����+D�:�݋���P02�3�-p�J���͗{��Z.�9�k��j��#p�2�-| �H��7�bcl��	.Ie�aP�mO�wE�c"�"g61l	^Q;_]l��161�ţ�@Hj�q��0^9ZL�M1���Y��K��@����.��� ��1����)��B'y���T�her�#��?Xo���ER3����f[NgIA1��s�I�4�J, N�z7�4����X�Oצ� G`��~�"�Bžt������Z%0]�B���`)I�<����J�,p�h�ZE�7��������J�F�뢜�" ,�I���/>���n��;RT$�%r�����`�0n�o�C�A���&�O6P��'3%��:�v"�2_��Թ�nC�}�"[1F "�I��j�)wnZt��V�x�bca�m�ɽ"��&�nOK����YLJH,��b�A+q��{�0��\zM)���J1;[v�h	[�3lg_13#K���>b�A|^�gL�֌�k�޸�cŏ_[{Rf�D�85�:�jdeg[�(XU��cK٢d�gY}�֣
�B�C^;b���a�q��gz��P��/�9�%��+|m�!����8$���	#�q|m0Y��~���4ϋ1t��H�I�Bu�7׵d�90���֊��3eڄkj��؛:���("j�9w��R�@.1�,�O<`��x�o����}6�|�9oٚ��u������.Bʸ!��|Z��p��-��ݤe����H��慢JfRn�o�ޗ�@�b�.��,W�z��T�'�m�6���c}�iI)���x��� �(Y�z*DLaq��7�@���8�dNy���I#䗚f	h"����b���mo�K��Ć`˻zv�Ȑ����SgeE��d�(�]�����;xgˋH���N�^�����*H�ų��[��Vj�\	;��{~&*�ټή� Z@��h�ЍV�s�[�h �(c��e�B&��[��:ıR���,�B7���H0�
j�GK�J�#P����Q0Y�vL�Ϳb�H��-ߡ�(6B�ܶ��kv��$�2�-�q4�vf���Ce&[^$���V:a���"��P�[u�}�j`��_}7Ҕ�5]�c��SCI|��5 =[�p�v�_�V3/��a)�Du�X�1�rk6��c\�b�`Y�c� ���fgMi���3�����mi���n�V&���LO��n������Ǳ�f`@N`�u�Qe����Z�@=o�*R
:[�)� �)��T�Qճ<���N`:����)a�t�ޘ����6��J
���o�����3f�ױ�GRd(:��) ��bbbz<5�`ʶj�V$����n+ ���z% �.�Ig?�P��2D���gy�Qf�����5�@��Ȥx[.��D���]�_�pJI/2�%7�x-H0*����y���<�o�s��u�4� �AJf&ż���r�F�k�#*'y��r-&�s��)�`��b�.��*bd�^-=u[Rj���L^��y��B�TI8�,L��iZ�ȫ륾&�C�(	Ch:���b�4���e	��-bb&a/;D�-��B�X�˘�o��!^�l;�ũ�(���e��� TᬈH&K^I0g5
Ja��<^����԰Ĝ��Q*�*6m���N]A2�֓X3�&p��h����DR!t��˝��L�����,I�,��J�#1�Qb��DC��h"���w�@�� ����]o2���/֋Q%�v�׵-�X�����F���	��������cX�J�0v_O�blN�9�݋z��sp&�3�٤ll�t��楻�7�\Ph/7���i@	a�t�D�K���'��Hct���R̷��I����a�k���2��6s������_~�m��2�#J�#]y�L�����u�JJ�������W�c��X�A��Y���H�_L��"&Y�5�4��r���h�B�37{R
�Z��5���6Ş�!�7����P����������^�g��^/Q��5�����@(�	mb�t��J�� ɍ���&:
�|��-�h!V�Rbut��I���7�s9S���b�G^���5�`˘s�\�j�NЗzO�u�GA"%�����`u�X�<�_)�#�f9�X,቟�U��(��y��(4�C2X��x��be{!�g�(6�J��Df�L�I�����x��&6�nZ��eb���oJ �T�i�T���x�Y�̶���/D/Ie���$n6��6f8���mD&fٍ(0�s~�33"2�����a�6K�;��f�+��.m�oj�o���ڈE���`��j�����E�o�v�[�lۭ.�Չ����� 8�"�2�ڋ$D��tڐ$�����i?�I0���h�c�L��q���5��QR@��ӑE��S<�b�|N�r�!-b߳�.s�K�!���h�->Hi󧒑-̺�@� �ˮ�Ib�4�2���RK�Sm���e&�DI�^*`��~��1&�I�ӵ�R�bMo��>�Q�Mq�(��&�Z�ms��K���g��ކ4��|߯��w� �2b��N��L��N�u���28rR�%�nb妛�%��8�;�f������	�5�![&<n?���!ptL���:B1D��}�ӄJ���6�{���$cy�_a���M!S(g�I���B��O92F/��^q^�m�by,�l>֍3za.�[Dͅ��z����X�x�7F,����I�6.M㘤"Q�f���Ix����\����f �^u��RdJE�b�1/~���BA�ʔ&$�̺�$��7����c
:�P�X�Gh��&&���'�FvӚ�d� ��8��J>b��lؘ��4�����V`������b"�i>�A�(g7�}iBXxb|Ql[��o��� ���J�w�7����Ǌi�~*m��N�('V��%܉�j@�� �Q7֚�X�бƛ�q[DZ߯�3�����5�P˔T&ޱFJR�pZT�:�M�t�Sca��m��T̤�Ab�a1��yo|�	X%�A�ɸG��v�i��P8��A��X+��������<_?�P7oF`��?�2����7� �A�Ⓔ�#�3y��	b�&�^�[M�NmG�E�kK})�x�oڤ��id�.9ֈ)��X�$���i4G ��IgS	!h
ܛt���A�1������=�����se�1�²�DlƂL6�0��Ɍ��$E !8�;��䗱Bf!�m�m�oQ�F���RH�(�.��� ľ�ًi�@�1,Ұx�Šo鮺Z�`�[K!$��f�&)�]��81f!a�i���s��:6��w�$ȋVa�f7T�8.^�%�5�k� ��ٛ������0�[�q�Q1�1��c;N�p�BQ9,�YE������[g��s�bY��aQ%F� ,ݑy4��a.��Ц���K�2���@`�[%b���m}���^�')��� �Y�#�� ��s-�� �N�L���?�bH�6�L�2�n��֢��ߵ��m��h3���\�WD��~�&�e���i��.��j�D)v�?viJ힔����g�Z+X��K�ְ���4����8�w���t��R�Ki� f�3bw��0�m1:�?�E<��_���L�}~�R�3����A`=	�<�*u�����2^`.�]{w�I)�2Y_���(_1)$����F/�(�x�����U��X5G��h���T���`*0b��vN�TәXd(�D�	�t�Ql.j�,j�-��J�Q,���5b&�bt�ս��'#=5c](Ke/��(���CۏzU{�:�7G�$�Hc��� �	�0�*���q#��P�5��U�iqH1
�b!T���h���"]�oi�JcB��[��1,B�������-5�eЉ��ƥВ P���ɖ(1��q�(.z����I��e,�o�ҍn�*%��n-4i2R��3�!P�.��O7�sQ�!ɉ���"�߬R�^�������3��ɧ� �X��)�0MQ6ސ�[x�����;g��A�KD���K%��5�9�-��:����';R���צ"�nq6uڋ��o�������G��j�x/|5e��a�1noZ��9��=�&jD[�9hff�8����9�ߊ[��3�i*����E�&9�~��$���O��/tσfc1���ZK.��zA�V�m�2�.3İ�6�(PXo��y4֐"`���v;�E1�`�/#i�D��m��d�p.�o53flM3&� 	��"g9S,�A(JN�'7����1�9��	lQe�n@��r�ȉYH��C7l
3�AIKx -��T���RD�Xf��gz	$���Y���I@�QZ�޶�p�ȑ4�No7ti)anm�i��}$�`n<�7��qR��4ԋgy��䌖9Yw��p##���s��N�0@�vn�oxH���yVqh��8�z��%ش��h��GVsl�.�Z�\%,� �,*�%	Phe`" jXKe��$))����u��J�����^�I0	1p7�S{�k�3�H� #$7Iv�ޞ�"Y�q&��B�9�o&�NF�~�0��A����R�B{>�3y�s� BX�������L^�G�b�;�A!�j�-�I���D�1��$1Z;�QhQN�ۦiۦ�����JT�`o�!���&T@�4�F��~u� ��/L����0Ii�����KRh�zK N�^͹�� t�n~t���n�\z[�u��Xi/���Rv'��,D���[�oo������LE��#�[wbA{�f� �*n��?�kRKfB�\�z�܉���Zg(��/��U�B2Cx���'U�1�ؾ�˭"�0_�<���K1qV`D�u:e�i��Hȇ��Sg+�׿K!�b�"HuŠ���iX�f,Ʌ\L���'p �����}�Oj�/)�~8�,`�&���N���T*	�`Mdt �P�8Oӭ�h$I)Q�C*';!��b�D���E�A��揳 Q	�^w��IL����[Δ�HX�0�Α����-���Dg*�t��Kk��]�㩊)� �I8	&�&*z�"܂P� ]KzX fR�1g4
 ++��ϮZ{�0�_J�:�Yo���4UTݺ�Xm�!"b�E��ޔ��s7����E`&fo�N��Bt"7��-��z$��g���"z\�ޯ.8ɏ�@t�{|�$�����2`l6}N�4���ǈ���+��ZqH��M���ndfVm��g���DH;�Pk���7�Z��:tޒH�*ѤzU惴����/�R�A�}T����ש�K{��J#6`�y�b'�C��(x'I~��|Ѐ�X6~��C��|m@ FI���zJ��.�h6��d�K��.L����H�Dk@��#v�jkǭD���yIC`��Qf�y�����1@�[���֖ �"���7!�i��RQ�m�+�jO	�'B{x�"�2d�Ǯ(xf	e�ִ�9��S�R3��o(B��C���l;�;��Z�dF�F/{�8���.	v=5&	�@� &��f�p��:�?Z�^��h瘶�ڔ������}��G��K�� ��P��]�3E)���;�:�pB�9W^#x֘`�%v�q��(������7k9dRaXYw�ӥ�UKȑm挘0����L��:L[��e�E0�%�]�ݼO$$	�U��e�LՁ�77��&bNx�Y6CA�f�G�aDZ�Ɨ�n������DJ�8ɻ�:�%97Is��FPr^�'N�E/CA~`3�g�0m<�~��I���~���,��F��j�\�8�_��*8��N����@]lx�Sr#	̎���/�f��1`��*`!o$�_�[�G3�,��8��JR'y /+v���Ő	˒6�-�Kd����R�i�Ls��C�ٱ���]4�+�"n4���cjHͱ���c���o�6�
f������0����o�X�D��?�3���;�bI�6�y;&��D���)���S�}k4$	Q&o�m8���6t��@�p����p?u�������ք���y�j�!6��ֳHǐT�u�8�
rL�I��1���i,l6�����5.�w`��RS�7���՚�[�r�PpeD��=,1��6��9�)�˓n���s���uw���$Z�m�� 2!qA3؈t�K�t/&���0�����u������}�P&`�L�H�pI%�h&ގH�ac��J�R�%�&t�49�&�L��DX&��b�"�<�.���y�'d�7�syɬE.Ap�5���-��p2i�ge��桩����0�qy
Y���փ7 Lh�b�bbzK��(���wޑfZ��.�%��3��ڂ��T�9fWL�E���c^zYj�Ő�:__�	�D�JW��Z�v�(�bb3�nX\fMGs>�L�g�#� ��Kc3�4ա$Պ"뗣�Z��c�q&y�������i��Kԉt� 6u�\֮�z!�gL�Xq��>0�/��1����`'��[�щ.���|M͋)�������� '�]��{����^i�g�ݺ�iW*���5o�/�5 ���� '�{z�, �N/��^��D�Yz؛o՚���]X����/e��R��;�����#?ʘ�7�Ӌ\��SFD�oiWPȴAМҤ1����v�0��׍rڃ��8����M��j��w:�/�(A�����i�oC�4K�2-��~*�؛�<��P�r������aw~�( �	6����bxT@	�ɏ�$( X��S�/D[�:�LJW���N��#���,m�9m}1I`BHVo��(DN]�/�7�$f�6{Ƈ�K�
$^���mz�%�W�����Cȭ����V�|���ۡ�=f~���b�k��F\�!�E-���C�6N��y�����ԼQ@�o�L�`4���o�-\G�~��k��J�b�乞�� ��7Վ�s�P.���G�]���7�/�i�M$`���3�yaL��+V�o0N��+�D���G�ir�f�X�t����M{�/cځ `����D��xu��-���^�����%1l��힝0`0)�V/�t�uV ���^�$���X�P�����2�x:�I�WR�`�\4�L�#��!���g)��N�j1(��;�z��ym�"�7����j���{E�H%+��6��vc����"w׵�F��>� +-�9�w��3�w�t���?sPE��ϬOj��1ק=i��Mz ��� ֹ��C8)0\���)����Q]=b�P��,��ϊua3���f�ʁi$A���'�+���q�v�����-��`�'�2��<M��D�����7
s=:�hڎ F�R�H%���r7���%��D.L��w������k4�E�����!ci��v�E���q�5�����|�� e��	2�j�3c�[�i֑UI����BC�!u/~<Q
����D�����a-�x��"D:A�ݭ'3@-��rJ��-�^�EB&��g��w��"&�Y�X��д�G2� F�n��}��}����L��9�i�9�?����7��}T^��SL��Ծu�>���!�k�ey5�M��|��9��$΋c�9�r��u٬�Ǥ���Ffͯ�4IIdo}��ڦ�Ny/�ը����	�>h%�1�s�S��u��hu!"_m5�Ss�<�E�f�����[
�ĶҖ��~�G������X@�ⓓ��ZRD/I��އ��\_�����j�ζ[��:Ԁ06�N�<bo,f�}�?�"��ݥ�F��/x���2��/6��8��o��bF��-�y���U��hKۚ
Ȕ[�{�.�p�ٚ�c���lx*�$BfG1�	7�D�i��H�V�qB$�F$�.�҄�B#�iH.aԴ�������;K2���*����P-�������9Ξ~��D�����GH�x����C���v$�4�ڔB�V���bv���
&!vC���J8�].�;�M�SY� ���r���ɹ�w��$�g\A��V�7��ӭ)Ci&ysJv��/����8�.K���ڥ%<^-r���K��R��$��Dm-]%�umHf��ک��2�r��"�d�7�h��/���v�C�מ ���j��-]+�}Y:���,�-vv�h�����~"���-ͱ>�o&����(CV8���*�,i�k�Y����隺`&=y�E��"�����u��.��jP��%���P�\����dX��jE��m���Ԥ#D�s�Y��s�;аr�l�&���K����AH�c5y��?
�����u�@@ׯ�t�6']�y�S�������qWS	��Ӥ��TIo1~�|QySm<q6�X&��E��b�jI�6��j$�"�y:kP
�Z|zڣ���&:^4��32�^�4�6�7n�t�5i�w��-��d%�vf��أAsG7A� 7�@3�������d.V'X�{ЀB@ ov��5&�B�#�B�s�QFf.�&��zݻ��`@���Lՠ�g��.F��7���JTA�"����D@�-n8�~�$D3��Oo�/@&fO����1y�O���m;�� 5"$�}hK`�7괪�4��D���6�2̾[T4 "@�( ��n�NLDK>�w���:_)� o���j��u��cE�Yc�hF$ƺ^�� (�F`�����vͣ�b{�_4��&���z���'��5�H�fsՋ'O�&�gM����sR�-��o})E M�g9�c�A��&o�D�:�gV|R+�Ϳ@G��3������5H��g��"�!/?4 �9�����F0�]:�n)W2p�ڕz����gj�i^����T+��}/GP����Z��n��&�{;S"ޒ(��g1�� �63��|����o?��9$�NǷ�8�`ZF?y�����{sѧ���g��W
�f��3�B!�'sc���^�7��oF���b��4� ���F�`�n��I�ZZ w�D���cO�ʮt^׋iIz!|��x�\e���Ʒ;U��ߧH���D��?�1�Z&�uT�9�o�|��AdY8�=�V�#P>k���[o��^!|:�C}����v7۩@0�M"���Q�����3�SOf0u6�H�Ι�@�Ӯ'ֱyb*�G3�o��N�a�d�#�c{x�],e����	��;:c�ԎoXI�LN�E�����c4�an��ݼR���-y�2P	�k�׊l豴�f"��=�J@�̷��Tˬ����f~��3���WN��s�@L�i�)h<���kZ�����(D��8��Ԍg�ޮ|���
@�~-m�Q>��J��Mo�={TX]�q3�ӈ_3���Օi����E�ix��hz�����#w��c�����m����Y��Z�:�����r��o�7'6ɵ�M��'<�5�y��������k��������-<Vn��"6����HP�^m�-� C��e� g�D1 137�~)zOY�X��ø��qN�/i����m����Fb�$f�j�~��3���ǵ�D�tt4�2A5��������)�>��$ۯ������RNbřӡ�zT,������2A0����J�<�����ugpw�ր"P��c�5%���3��1z�am�t�f�.نi����*%Q�3��7��#��*�$Ύ��͙�� l3�[�tz��C:N}�s �}�����e��w��L����mE^�F�ޤXQ����H�F�����M�z���HlDZS�(]�1�QfM����-���E��Ǌ=O{�Ia�2�,N^i!���3���#k�3��H��l��ޒ�4��]�T�s�{S���L_�@Y�Sn]hB��Yp�ֱ ;����$��o;T�=t���NH��-�'�{�(�ߗm�kP̊fo�X��4����X�l��.]�LkMN!{��@vA�u׼R�<A7�*���16�A��0b���kKd���%�̤k�E����^�7*@}?�
�$ �-J2m������.�t-JЃ F�Y����_�Q�Q$�/���HD��ڔ��o8����E��X*4�"��<w�H��}��g:�}t跣ȯ�4���x��������Z$�7�H����*�-��ƻ�ژ�nC]�a5�~'n�ttu8�P��7���t;Gv��V-�]6�^	�w��O֫����\�L뉏<M*�1ý,E�o$�ԡ]�Zb�lL�Ʋ��}�d��0y�:��=� �W�9�sN�!��](���A߭�f#�j�X>/�;���*�p&O��j�MD^���f���MI�ts��h�����`���qh�<�撒�u��4���&6�։nc6���i�k�z�E�"���[/�|z��4�!����R���b��o:�zN�D�d��I1)��>��d|���a� �/ko���r%~��%�m���rΜ�n͵1PB7Ky=Z�Ē��0�b�{:c�;� ��6=}�-�t��j�a�{o�A{m怓y�-�y���fڻ��sp�m����
2Zs��h� 3���(�M�=!�S���"��q�l@��:��I���$�>�ԔO�j�K��=#��R�%2�s�u)YCV�z�L����O�=�Sss�특
6/��,���Ш�i����E���բf�.����Q����g;a��.K�lo3��`��Bm/ֽ��ĘӼ�u�/�\F';�=�H�9�w��$���O�(�N�ZM�v�3��f';��D&�c�^ P�Ւ��Gb�Y�sJ������t)-B��hZ6��5]㮳�B"I�:�J/��}��F�-����g�(���u�j3'+m(���M C��{Ԣ1?7ޠ0Me�q>?M!7	�&`�|tg��_{o���h���D��f��\ ���jS��k֭k���qQ&_=�ir.���wa��*�X�������e:͵�y�֬�%7�5ԃ�4�K7��"�u��"���=qPm�Q%�r<6����I9��ݨ���f-�!��`��nҸ�l��{�;S��bs��jU]K�S�̮�n����F�5���o�\8ؚ�z:�T���N�8t�4�]~���$E����ED������+����*@<˟�Sg�R	:��p���Ԑ4_xOZ�7�v� \yo�4��z�pb�fgr�h@��V�:�7�r=R�k�,��j����Ǵ�ɡ��ש���6C���hu�C3��ށf��3h��n�NՃ��LDC��i�֨�cL�;Ա����yлءF��8�9�Affb'T��qc��.܉��g-~�κQ�#Y�[������=i���sc��Q�~Ɣ5[g�F�3�3M� ����y��Ojp-���h�e�������پ[I�b�:���5y0<e�m�  R-ε'B'<��H�� b�9�4�#������ �ڈ2ݱl�t�1��l����Dz��s|c3Q����m�����,�zLڦA�,LN���L��X�o��hzY� Jx0[\� �Z����0J��F$�o"
0!�g�jHL�s�����ּ�Y��Ǚ_��\�f5;�h���H��� �R�y���8�/cM��{T��,��j�0g�l���nA���:���)2BCf^��h�L�{4]uML���L�;ǧJ��f�(H.����飦* �2ש�u��0r�ؿ��0[���Q�������7��&��ٷϧ��1�K���ؿf�"-��!bSm綻�A�6�sk�^��Qĳ�hǥ`���ڔ`#$�q��׍av�^e�K�3�<ЀE�&�j��#D�y�ϧ�J�U:��#g��}��ܞ�3�   %�=\��k��}�)L�1��
����D��ų8��� ]�N!�fuK��R&X��J�F�gE�Phm�_�
&��o�}3�N :gW~Z ��Y֥��Dy��d;J}ʜ�������4"���*W3�4;�=Y�ZYt:PS0kҤ
�9�JB$!���[�� ����N�"mF��ӫ��#L�����]%���?��J'h�hN��EU��;�vڣ,3(��Jj�]��K�9�r)��J��C����:�uU����U���K��nu�Q�����H�D[��G�R	8���8�Ց����*x��JȇG����a�g�?�#:v� y��sOA{q{Z�%Żm\��Hck�T���b��@��o������#��d�X^8\[��iL��M�t�$S�;��4FE�}�{��u33B�ih�BVv|\�@�s��	ؚ@b-�}9����N�֌$\�O���s'�y(Yf�H�9��
bmθ��7���c#���X:��a"����`�3�ԑ2Y��x���[s��i��� 4�bMg�Ԩ��<���PJ�`�̛Q�&}_�T&/VQ�`�1���+��L��k��v�,{y�x�SƏEd�c��)�`�Z�������[￥���K�'�gV����Bv3��c~���N�!���b��Zs��~�+����jK�������F/��F$�gx�����St^pLS��'0c��.�T<��ލB�/!�<v�5�(�3��J*�U��EɅ&g0��ɨ	2�߾��n�VQ���bxդ���{� *!�7us�YP�������C��� ��O_50ģ(�b�֍�1`��% Dqť�]�T9��a�L�8J�9�smy�Zbh]�b�1�ŪQev��-|�Mͪ��rk�רWB�)r�Ҥ����I�1R	$�#��6���iټ���Rp"'I4�R�˛��&&f-��R(Ś���G�4�B���H&I�>�1�� ��j��7��sQ�fgi�o�@�P^�-o5
Ǧ���-�5���GL�Te�Yn�\zt�BH�oEb[ϣ�\��p��u�q��(�2ݻ��	jdaf9��ȹ��LQ�ng⑆Ƙ�3m1Ar`��1�L-ٶG��E��"�q�?w�6�����X�Dl���x��,�S��F�S\	�N5�-7�`�+����M�q��X���\?η�X"bt���5�b I@��ӎ�����0����Z	��+����q�#__D1��	$�����A�U8ni��QY �X�׾�� :��c.�\�Ý5��
ES
�1=i��'p/�f��7�b~1�,�M���Qr_>��j�E�,6s�qoJlc�,��^?�:��j.��Є>�臫���m:�������LU�K,���z-�)��Vٮ����( � ��;�Fy������ط�$n?�"L��cٚZ����-�o~�×1�SZ��q��"V����Rb�}:��H̚�J��A��~�H_{�zއǖ �Q%����7I�a����4�� )��=zR�'�j1;�ޱyb* '��]�� ��5ԥ�����F��t�7.�oׇc�Ғștm�`�8ə�2#;��3�(Ct��Qd��cޘy�m��~{Ӵ����1���&smt��Y��gڟÊ�
��oE&�	rkI�x�@�w$�{T�H=MNO����?�/�s���X)�K�0��ę�AY^ny�h�z*�LM�	��Cq0%�ϏZ��=/���*Q�Y�Կ'\Z� pD��iW
$s��$^"��r�tc�?f��1w�ZiF{^>5źѱA��ut�?���؋M����L�r��ޑ@�"'I;y�k&C~綃ҵ�fb�G���0ҀBR�HǊR�q�4����z���_]���X5���k�B�:[��阈&w�~ia7��)s��@a��!(g��� 1�bv����b9��윭"�FÛcg���3��bfo��Ox�M�5 #|q��qoZ�|ָ�E��{��T��н�V޴�c�O��`�����[�p�K`@�!���fv3?�puN��hP%˿��-�}oҀ,n�3B��[X1Jq6���I�|/�zb!�����g30���4ޱfo���k3��($I��� 7�Pc3m1H���g^�-����X�$��Є���~�^��f1{��鍩���K5�nG\��-"��>*]�4H��D�ןym0�x��и$�L�k�>�v9*����ޢ hz�3�3Jw��6t'�M��q�4L���:q���� `���8��d�]N����/2ou>(�2u̓�����4w�(F�gw�1� z���L���l� �/H�H�� uޠ?-���v�&t.��b%����/�ud���*���٤�y{^���sγ�s|�׽���&P��oh��JuGI��1�c[��R'�։�'1�!f-���z!a|N�G�Պ�l��r�V�[JD�˴�^se\�O�b�;�θ���Z��D~�10��T���B��k�!��{u��Z�L�58�_�Vq/Y�'z2=:�*f���ڍ�E����A���A���LTx��� ��f'��jI'�:b-vi��P��Sl&�.��s;]����y߂����LRĒxg��֝cϫk���<)�G�אE�~�㚑X%����EI2���֢�fq�-�F��m�n��|��Fw���� ��9��|�L��{�2l�a�/�R�Y7DM�o|��*����t�km�������	ۦ�O��J��u^�p��BO�������Rd�"ٽ�����ӊe���^�4��4���xs�*���.,ފ��eYu0M�iW�ϙΖ�i�)���L�B^HT��O���A$�1������ԩ)?ȩL��n՝�Z2^8{T#�}��^�`��7�X��H���й�M��l���[�j�l�oߵ ĝ-�I�my�m���4�f؋�b��f5�������:Dq4��/^��AX��ԊnMn�$K�GY�څ�?9�Io�����6	Jd$��v<^[�o����O��mC#^q�C%)���Bs3�� �&#Zi�>�6��4$�OF�I(�x�ژ	]3���|�Q����f��-�gY��o����)3/^fi�s�؃ަb���� ٙށ��;�������\�]��4��wd�T B�|5�kQv.F��$�ў�BV�!���놓0�de�(��#�J���!1}k��3�C��zxH�-� #1��*آ0f�-�x�JQ��_�v����)����&�َ�7��h$D^�6���<y��r<�F�9�������ID�I���k�g��
�2��F_�͠�K8�E�scO���� �&�o:���=�ĺ�)����� ~�1����Q(�6���jD���ojg�؎=w�$m/wk��*���q�i"�O�D&oI4���Mn��}��1ݢ�m��4b/��49�G��3������y��<��n�-\�;��42��T�js�W�bz�'���������9��ҙ3�9�����(%�����m�� A��/nV��6�R�4��9��4�����J@�s����P��=foH#Q�M�Kf��;�����Fqxɭ�G����$���<�"��&'F^]X�u�r�7iζ"�����X��H+D���>hv�5�j&� 2�x�\R������S;n�(,���/髮h�Ou���mh�$�!WKm�F����g� a���lx���/�i�-�z�E"ql�K9����>iJhDu�;�R�X1ln��B�B�!|��K�B� IAd�E{�M��K*ڬ�w�<����ݍ�?䐼z=�@�'��ǚ�8���=5�K,v<U�a#3�@����*tYw[��U��4g�#- Cm�#�M(X���D(ZrM��J5#��(�39r���nw}H*J �8g)?�@���K�Y� ��̓��JI�隅��_=i�>Jh&Yg��U��5�S�ؓDpE^u�Z N���Z�ǭ.B���Ҙ��c�I��aJ�w��1�������.b&��j2"�'K3��┶a�/h��ڲ,Tam��.L��(b�����.��X�	�������P"�E�����	،�2����'�zT�s�}����g��$���Í3DB�21 Z|�,-bLE3/��P�;�R���v"w�]�������T�,�oס�N�Mft7�5 ����x����30-D��m�]���"���Ƕ�&!M`Ƴ9~�Q�!�f%�B�!Vr���W�2�sZ���3�Ƶ)�t|��� "O��'���ϽJv3���ڔ8��Wd#�v��&'V`Ͳ}Qk\��J��y� >�Pb-����eto�Ξ�K�\���8_}�d/���4Z6Em�����HD��
%� =k	N�9Ζ�Qg��զ;�����-��%�x�
@�A�K=#J0��ÿ�ǚ,
ɉz��R��N94�;�=(�P��|�����O
��`Yl��Ɉ���jI��X�?`�z�=�X��Lw������H7S��j'X�??��9�U�ng\~ޙn��qQ�.g�D�/����?=���еfV�b}��܈}1��y�������1pv���m:c�� �m�����(��k�H�1�)Hi������'�k[�^Tb؆��O��N8���DL��PY����o}��o,��-� vtn��K��x�멾�t�_��i��bu�ם<�t4�,�s|�v��[j"�)��m)\�������+�-���5.#,J���m)E&Ƅ�|�ʪ���,G��!L�Pxe|,�8��D�7�ŨŅ�!,�X����o&$�#n�f K +��[���ym3.��֌���3��g���[OJEbŵ܏ϭ8��w�A
1�6��P��5/�sݚJ���KւV!��Nյ����&�7�ϥ�F�qG���x�	��o��Qx'���b#2���W�r����N�3h������]b����K7�?��(6e�(ğ��]������3���iPw�I��Җl/�fsހ��M�������41	NH�c�$HvޑWx���'Ҕ���tޥ(F�@�7�jP`���W8lkI1t�i�fMu��ڝY3kkx���<|���7���M&D�qgJS�_��Qgs&��衸�!�J4xgog�a�������5�QMО���Z�
f׼��ִ&�cj%٘�g�bhs82E����4[���LZ��\����i=�Vo������	"�O{���@2����x��]L���EX��lO���^crs��Z���3~<}P!O;��{�t�"p��cGja9�8r��J��k��Z��R��X�� Z��� _e.ߣ�/i�Do���F��[9��F��:��0�NN�h�g8i�3�[1�Hb��7B��sS���;Q�^��|mW�s�@��M�O�"u[^�ue:�.�_�Hn���FA��PD���Ιڄ��fN���#��oDF��κߊ�b~qϥ$&���Jd�]qL-�|����y����,Ĕ���:�Gzr�3����]}�\������Pbm��(�Ͷ���Y��g���:'8t��M�5�~4���)��|� 5�n�c�N���R �,�6���7��Z&b5�:�Gw���LFn��������X��}�����(	�q1>��K����;�>�y�����x�ތ�!Nz�HMR�0�Ƶ$7��X�Sk��L��'����D�L����J;�:��� ݤ[>?z�������4��މ���ֵM]9�H�{��[��N,A�'�̝i����͵ߒ����oBU�2m��� �I��Yݽ�z��X�Z�y�`�=�X����Ғ�7��{m�Rݒ���u�RC}��R
�N���b
�O@��H���'9z���A�b2_^�S5kh�boRX�u�f�
�3{�}3Chn���F�	fٞi$�9�s	ސh��X�m�a�Z|=j@��m4(�1����2u��Q�ש�j�f����R^��١[���r�D�#�]��)�q?�L`&�����?k�  ��P`Ds�٤R��ُJbPY&��z�4�FbiRK��8ڄݾ���4]l3��z� ���-`����PÆ��:R��_7��4�J X�u�fs�S"$�����ʜ��N��R�[g��oW҈!\߬{�ʾ_�v�d�%��%�;?��r[L����dE�mk�!���c���dT:�;c1�5R�^�	%DCgU���;.�J�ډ,Ix[��oG�z��@��[g���/u�/;�Ǌ�hn�QI͙_k� �e2'��R��"z��m3Hihm1�%P��C�?M�lA�^(D�6��Yq��S�Ҟ�G��&iC��}�8�� .2��$�>�.ёбnW�M��J�1:��<�]���̓�R��)D[z�q���$��f'@�n����JR�7��԰�o-������:��0I���jXi��3%dm�x��-@��\�5
&/���@L���ڠ؞��V��,�-3^�&�ownz�L+`���Se4=pޢü��n�mCf��qS&�[�_wǙ!��y҄�p�;�:w�4�f׬.Ţ�3�����s�Y���hSA��<u�׮�$�D�42�2G��@Ҳ]��
%k<�N��V�s��I)�뭨@M�6�4	D�z�t����8�F��f�XǑ?	��`�|��q�3�h=I� ���+LD��zF7�H�9� �o!{f7����ו���h��^�']o�AX��f^�`Ҧ�׊K�q.�x�n�B��-����օ<�$$��� f� �����P0)�"�#��-JF��Q�7�v��l��z�g<٩P�ϥ�����ǿZ:�N�ܒ�؊�n"i{��� �B����PdͶ��Ka��3zl"�ŧmf������ � DʧZ	�3�EbB�l�X��(-����K�d�o�^RE��"T�x�
�6�Df��|/�H!7���|Z]ҝ0i���fήd�歈�qm��E�u>	��!v� �M��)km�қ3ow���K�c:����8��>���x��o��Оg�H/��Z�w�W
���,��F�����)`�b����K#vy;��Ed$����~���o�ՎԥHTd�Kw� i;����
���x��)�T��~4�@n���4�H�a�=w�(4�����t��Vg7ڠI����ڮCVv��ځ�f��z��	�����6s�Q� ����j&m|lT��٤n~���D����Db�hd%�E#9�ך.pb;o�4�U��E����W�VZ���M*WB��;Zo3_�S!a���ɦ�ж�m����L���D��M���䖆}	ם�S.ɼ�����b���� �N�q�%;xlf��E�X�o�b���mΑ���Q����Y"&�H�8�	�k�Z�:Z@��⋚�ӬP�~>�D���H���_3�5�V��.���w}��w�Vf;ο��Ez4J�lF�^w�J	w�ڃf}Lu���j��D�oR.���*��E\'Y�GV�!bO��(v�����$؈��֫�F���e��~߷������J����K1yݱ���`���}{M�i!�K���ST�NLmS��A��N����~��������*fg7'�a�X��cv�[u}v��-D��v��g�V`��~�?��r��D�oL0w�X��� ��~̴�;�!��R�XĽg��(A�o�X	��@L_�3� '���E1����%1��=�N$I��Γ��1�[DL���cM��Pk��T�lk9�o��L���5H-�*�yD�ޗ���F:�J+PI��ߴ����f>����z��	��bfh���˫�-ަP�7�C����	0]6��&�k�ұ ������޲�:�͹�'���G��I�������<vƱ4�J���6�BQ���!�`��R��4���go�^�#3�� �-o�zR���ޗ2��ނ6�{��b�o�w��H9��̻-�qԩ,�O� �x�wh&�H��8��*����d�ш�N�@�����;oM�"v�����o��z��1�kf����1��Ib�L�l���x?�`��e�Ͽ�\Ƴ�]yi�����!b�ƽJ,����zT�$�d��Q��7�moSi��_�$M��ҝA��FY�G;�2;y�J����� �4[�sx׋^�nooG�.E�	ſ�����l���������$T$19�/�ڊ;!.𴴲W�b�:g)���x��K��j�n�4�l�1�q�I�̺t`D�Y�>��[�P�\�с!�L����t���q~���X���=w��jۺ�H��F#��b�����P3��q1���3�7u�;=��p�':�����G�4��+1z����m���������ӯI:S`�ϼt�&��y�34�M�bq���A���[���b~�(��6����>�_�z,p��Nq}��L����١�!���8ޡp/�# cmu�N�_ء��6�J1#�����N� �������Ґ��|� ݙ�j���˴z�)g����N`�oM<�]w�DQ�=�7or����ٴ��#�v��6`�����w��,�Ngn�b=r�D��f#N�CR}3�#O�J'�\���m�%��D ��}{�U���ܷnj��m:�4Y�����3����m�"����� X�K���F�I��N�](���z��=���-����(���NӜ��T��ؗ�͝�� `���{DE��H,d��F�2��/;}U�Y�� 1�#2Uݤ{MK�榡1��^�$�`�A~�qLM���~sm}0����V"L�ah 3b���H3�cnL�ɛ�G��=(�
��d�("��L���"#<�N�w�]ܕ�Y+M��U��*0Λ���������N���km��ik$G�B�.����e��ߝ���ycgO�"+˼��\D�fm	�V��/����1��M�w��$ H���7dq1BK/h��T��3��o����D��� $�vS9���7&cSZIF���5)�B�u�bSk��E� �-9��z�������� �<Q#sKJ��K����8z$�9M� ̧�O�j� �N1~ӆ�DL��g:�L�Nb<ڃL�ďc�3@��{8��H��=�����CR�e�q�ǥ
ؘ�p)R�`��[�E��1�6�-  A����%�ts��. 8�%�>��ʤE���w�N/QL'u����b)`���O�Y���"�,���ݣ	Z�t����iW:�8f&�J�3����z�:�3�u���B$,�.^jr_�� f�*��Ǘ�� �QWfW�����D����KЦW��9������׵�աkI�Q�D���I�%�|e�6�����'^~iH�;z����1Ad7��4D�ۜ(��>�����ʐg���;�oMShw�m�@BMfg_����� ��2���I2Β�R�1��uۍ��!YA�D�`��N����!<�L��w�&;q�zL3��0��ܯ;�%牉�c1R5~J&C�8�B��yأ���w�K�����1��������ڱ~ՠ*O���"݄�;�朚��6��4��Kf����g��x���!��w��O�.5�3��Bɿ�Z�|�޲=Ooz ��oi�U��)-�x�I����R��zm#\��h�L�3�8��\~�A�����4B"/!s��LOc��c*�ՠ%C�j�Ӗ�D��ȝy�=��Dè"b]1�.�,����/)d�o��~�X��\��K�3��ɂ61vޚ����F�}9�2Q�����D#KY/�[���3n�h#w�j%���[{oF���M��$$nFj{� :Q`n�g-h�8���|�
"m�\��b]��@A�_��4�4�kP'p⡇_�h[Fb{���^'�JO�>�(���4����-��+D=��ҲTJ������Jq<��=��C+�bϟ֨Ii7�\i�)f���;�Pc���0 #b�ҁ��Y���.$e$�m��-}�R	�{��P,��lG4�<�3��f���>ߊ�d	�����o�R1m�D��"L�wJWu;��x�L�ʷ���hrжh�A&�>(�C8��D�szc��z�h*^�~��N����Mv�jDfO�/�M���2���5��t��� 5 �����_ؠIP��qڢ�BMz|]��H�k|�A+�&�{��bB(��C�Q�*"0���P����w��Zy�sփ������ҚS���=)�Xl��1�+�[��՗ILI{��A������(��'�q�4����ö �_��-�����{qK%��Ӎ(\���XIN���)��߮�	"ͦm�f���.��̱1m��*Pc��N�1��[�>��;���C X����Ε�����&�b"o�a�'�ڋ�=�w�7B�h���c��X���s���"�d�}�#fS��w4�m�k$�̮�m�f&t��3-0	��y����I��N5֒my�W�9��c�;R��m�%Lw/;�S`F��g�z��v���]w�O���:Д?b�7���q/�h*C��������� [�m�v�Z/�Z��,P	# -�PI�hLv	��=:�o�:.Ȟu��@S�Xδ�{mB1�����	x�;�nk'G���~��ːNczQ�s��D�mJ,�1����Z�5˼�(fb/�ܞz$JKM�r�
N����r����
򩴾�� ���~�H:F�{s٥5yE�� 9�M�~�Y�9���`��Huڍ��/�Z�"�?�z�e辳��5��h-7��sy�*���'A�@�7��-��@�go��Jˉ0;}/:�:�hid�',ǧ9� Q�OL��5X-%�j��;␁ٗޅ��8��Ь̑}cCm��!fo�?�%�/��jF�_�q�\BA�4�zճۿ��Z�׭:�!��z�88��b���`��|�"�m8�u���j�Q�3<�h�'�ǘ�`�&�����"
	���-Q"2O�r����~�2/�w#=�� ������ 0�y��� �'7u��R��h��4�� ��Ks�õ����`#��od���� � t��l/��m��4AI<���qc�!��H2���VzE)Ჹ�4A�dĳ�����uS�����h�fX���0�Fe�DM����a$]4���s�Dy� �V�t'֬�L���ѩ\er9㝯�"�io&����-�͸⌈I�~�-r��ķ	gT����̺��X�GX�U�v�K�#b���J����v$��W�kS ��[ů�R8q�B���&�M7C�?�(�Y��̘�EN�:�xڈst���[,���%�M�:�3��(�� ��Oh����DO-����1��gj����┺Ɠ@m��t��&b#~�7�at��i^͝��E�%��9�����BC����~����m���W��M*��s����;q�J@��mtӬަXuCm��/�) �sjUlL��v��]#>e���c���n����ݙ��_�7��4$���\�Q3��c�V���+����3;P�gx�]�(PP<Fcj�H	�ߝi@-�%ӿ� E�gL�O�H��[��m�ͣ�l�5xlQ(��f/��D�M�^k)�fg���6nQ��	��JG�����3�4Jk�I �:Aq�G�+3�b1���hd�ޥG�b�P"�h�Y���nZ�A�bϦ��w��[8����j�~��Xf����h���iS_$�[��x�Ł+�ŧڂ�$�I�MmC��U�Y��S@���q�ks�b�B�������֝Wo}���Wwa����n���u����$�pX�O�H�$��*�����O����2��j����zR,X9[_�f��X�ɏ�M7;�x��Hb��0�u޹	���H��4,�"q��hz�ԠL��&-~�hK ��mD�����Yr�8�JAKi����zѾXƮ��ӛю֩�X��z�!�-��H��c�Br:[�H��/���Ќ� �A}D-Ф%��Z|w��<���
m��I�ͱ�?�]���f�y�#-�Gm�}�)uY��� H^o�{Sl���֎�Jf;xއe:C���@�&,!~^��6�cژ&�,��zI1r��N�<з�i}qojl��r�ED�Jp/��Ff�fo��D�2XB$Ǜw�����u��[FIL��|F����Y��ӭ��p7b{i�A�,M�[f��XW�<o�A�$\1�xj0��1w�}��;��D�ץ@ټ�/��*e�&X��w.��g m%��#gh����J�o|b��EW�ʹ��A�����`�/IH�)=#^�7�%J/����QP��[e��v�Bd&!�]/7��g�-��b�9@t���+����,��÷OJ���z��m3��81����B+K�D2��]��oؓ�C$�!�1⌥�m���E�rd&��[�Yy�ޥ�F%��o4t�G�Wz	9;�L��]�:���Sˈ���D�����$�g�"�<1ζ�������ntc�b�������00��U�M�w��X�Y�D���C!sO:5+ua��>����$��i�X�����Gl� ���ډ1��{եy��?�2֬/X�<G.7�!m�u���I�}(�8|Zt��6��z�-��-����O���Q��ڥ���־�E*O^Ry���D����� (��g�߻��7�eKo��*o��ׅ�jk�m9�a�֠0���gM���:�c�*� ��J��#��-RC�~��76��s�Cʆ��u� �F������۬���_�������j�D��.�"s���Z������"��4x�:ѭAw&�~'���c9�zSb���11YU�4?5<0�
HՒ��j���n�o���B�/���4�����/��P;7�|T] ����Z� �mq?��V}n}L����[�/*tb�����k��D-����\��M����ǲz�mP���ǀ�$��"K��@��u�iY����E�W3P�p�I$bn�8�����l��~&�&ͭ>
M��;��#4c/y��X����PE�X��'żRX�g���Y�fn�mJv#��}�BE��n�P���s;�9�Hi秮h�u�3�L�����@�<TFl_^�=������un����`�1�Q��r��M�n��q<��j�%��y�������ޘLCX���kQ��2���o��7A��^��M����~؁  1�^��M����ޕi�L�y6�Ӏ��r���Z�3�����^��<%�av`� 1I���>�^�<Ș�-1�Z����,,{�镾[tM�D%���7�_S�Ma��{����	u�����/�������$��.�y�&���z(�~}|2������e�ϩ��:kM=�*����P^��R��R�5��)Gq<e�P!�\X�;���1������u��ՂKq��)C�<1���@��8�!6��ӵ(:�wK�Ж�#���4 ��j,_&u��Dmo���MӉ�33��=;�=i	38�1�����0.�s�A�9��j`Yl���8���u��|߭�GT� ��J���h��!���oj��8��?���O��PF�B����H����1��O� D�����o�T4�~�XI�φ)��aͼSb/��k}�$__]c6զ���yh%3h����;��zYf�d������(O�f3ͨ�4����.M�3�'�Z����J';o���Ǘ�^%d���a
f���q��K
�3����+�g��馔��02@ܟ^�l�"w�I�^zղ�,�ߵL ���PQȤ�q��b�2�@����4���tY����R�MW�c���Jf�*s��A�m���X�!����]��2-�i��r߳H�[M��Z	��s��W �E��_q��&����{P�$M�Mt�RZ).dL9Sd5�Ve��� (�#�]�����fw���[��o?Ϳ�&fu����x9���A2Z�i�Z3F��"t�8�͞�	�[G���-��إ\�ք�v��� ��~k�Z��H�,ɷZP9�T]���ix��AgZ���Kߵ
"Lc���,�������\QE\�v���Jp�m�P˼Gmq�D)I��O���Yд:b�"Ʀ�F=k!�P��]�������=��b�� ݄�s��l]���ͺ���^٢0�Лx'�z2����N<}Vc�ݼi��׼7M7��"j����Gtr��O�(�rXs>o�8� � ��ǥ .�y���|��4'>i�de�]]���(��W_����������y:�Ҭ3c�>�9á�m͵睻P�H7�9x��Yf��clg�I\Al^oiӊgި�z�g��FI��)���k1���\c��<LQ�nk9�_6ҍ��N���0�'mz-�7�I��lL{P�S��g�=�̣ή-��(��bv1�L�8�5�Z��t����m��zB�����r�M�ԁ���40����s=��� �.Ƴ�3֥&;�s0G��)�ʸ�z�\���K�����'/Ym�� r���&D�� a�Iﮙ��x홽.R/�Mt��J]$�7�C"nz��%m�ݍ/��At�Ql�^?ZB�Wf��i�h��9�J"��!�b ��%�=��A�2����I�K9��[ͱW��[JjKI����#�_IjI�����E�N��-QI��1�b�5,�BS�����R-�^|{t��BRo�zo�YZ��؏�Z*�NҒ��g�D.��{��.qm6��D�_�5��F��e�_��X\6��đa�gn�p͌o�X	�뭦#��!c�6������Z���ގ0-��g���B, kh����i�$�3/�3�5�� ��0* "3a�m;�K�˓�p�*,F����6F��U�D��ïo@X����P�Ĝ�~�	�'}j�!%&����d��j"���إt[��J�&����d��+�X�t��-���ǝ��?	��>u�j��qRܕg���Kk�X֥��5�z��.,2���(^_�z��)$�)r�8񚄉!{�-f�n��,O��\�x��L�Oq�Y��X������ٹAw��}�z�K#6e��֖���7_#i�g^���5;|հ�&�v◒��8�oB H1;?qB��L�1�~��?�
�Cf�o��E�[J[&�����C�8����M1�#wF[cH-��R�/�4{>�Y���J.q)Z���^���0['�� =���,=v���0�"aQ�w�i�"�X%�n=�kZ�-���@��ob���%vy���HfV#$:�ڂ�Γq���!��n��IA��@:�Z����d����m���$4�[o�1Va�	��{}̑�>~�Q��P���{���&����"�h�HA5��oZR���w)�"�.�^�S�mF!MQ�:���N�O�9D��[L�I�ۦ�Z������|>��5k�c�h�J�V#�|�\v�Z��❳>�h�N �&�R��=������qP��a'^�F����"�2Ќ����������6<~{T%��:S�}���%،\���_�z���ыTv�gmZ{1���R�i1����+9�� �3?��G=i@����i�:���IY3>׎'N�+��ݥݜ���P��3�6����T�"�f��T���d�f�D��jA����Z�ȄZO���R�I֔N�䏧�9<��Ff����峽@ȉ�mv�_h\L��[��g�xzYۡR�K?��׵A@��iq��>�a,l'.w�����bX��P�ĳ;;8���9���~�+"����B&�cl�c�l��6�i�������*L���ͪ�"��3A�Qռu4h"�Lěo�A����ؽ鼣��qHH�������du� hPIL�^�XN�GO�jL^']�@)6)���i1�\�a�:Gi�RD>W��O��d���������'ΙަX	��:�����׬�bt�[��P�L�[9[��j���i{��$�cP"�g�x35t\t�X��qf��B �TAu/l�{o1V�t�SE�;i}�W��>q��e���Q����!�a6a~⁆�4^�{�J�Ᏺ�\Oa�ެ%�n=�h�G^i���w��j2��'�s�	���6#l~�)"	�ԑ ��קO�WQ���J��:�(U�괁	.��zt���<k�h-]��b3o8E�R�)���|�pV6���� ��>4���4��P�Y�:�^����\Ν]�=��ȹ9�:�<u���%�(X'd�6<�)�|��r�̝<sH�-�!��4K����0S�!����HRIr[�ڂ[r�J�̈�ro���G>�q3_�J6�o�jFZ��j���&B��C�5�����ڃ6������|աk:�ށk��E��]m47��ڤ�rU��%�o��Ǯ��P�:z�S7:=�Sp�����*��Q��v�H���q��梯���u�K_ژ7~��5p����Jp�tz�� 4���"�#�Ԇem���jO轴�@$�����)"�8�� 3V���r�����J\���I8��Z�����zTY���ړ&��æ��+x��{y(�}�����U���Ҕlj��[Z�)p���D&�}��k����2ϖ(M��:��*����5�� jy����j
���/��R(����D�* ��z���a�\�ǯt�ɓRGK�چ� u��s��,ͣ�ݺR��mU7M������7�jh�)���E`�Ӝ��,��(`�;t���ݕ7��x�t��'^z�bCm�x��j
�<�v�gQg�8?T �[[OoP�$&uh�Z3�m� /���Fa��z|���[~�A��0��kt������r�&���e��3uc����W*�Z��4HIԎ�w��k;��@�sr� Jxs�ݫY1��"_V���pմ�u[x��J�cX0�c�n�Ж	�LΓҤTӺ�mD����ijY��ޙs���g�j.Cv,���ETƬ������?5!���H)x�լ뾾i%I�ޠ�����V�ѭ�c�zT���OSΔ�2��U��lT�nOko4���QKg�?��	��kNh ̸�sEq}y4������nm�x�F$y���SQ��WOZm�����^��[ۧJ��&vr�U �[I��!v'�@`Bo.�iP���\����sōm�(����}��$�xI	�9<��V)�r������<'K�����ХA�i����&��������J��#�ŦqQ�gx�����~����t�h�Ke-�T2��c���#�=)½И�K��b�� !Y�b���sQ^Ï�� �f����o�E�����F�ϥQ7ޤ;�O,����o7O��ֈ[��4�.o�x�@[����`Y���Z��ƾ�j�|oe�7��0g�}����ǵ8��u��i?9��-3�tޅ2��%x��N[#�LO�T��Ь/F4̴�5L�1;Z�S\[�tޒ�{��^
\^#{�%�u���Ѝ���Y��_٬s?�ܦGrі*Z뉧���&\{R�b��Yb�8�b�{��j�c}*@o3�f�3�J�%y���t�Co� �h��<t�Ӯ՚t��Z�M3�x���Z7�u�gǥ	Y�C����8�١)&}}hS��8�m�Inqş��@��b�|[JL�/i$֋���}����o���������5����d+����ٮ�7���u��n�;� 0@Ͽ+	��o׬�o_h�^D�.�5(���,�3w~��֔�/�������Nl�'�3Xk�g��Crf[oօ��3;����
ʮ�gM)Є���iϓ�0�P���t��W� �����S� cby[����,�1���P̛e�3v�_zX�BnE���۳e�� �h��T볛��Ojb�-y��I!b�ZH K7LG��ҥ�L��m_:7�n("�N��뚾��e�I6�6럪av���F�dszP�/ڢa"3Yt��iAt��Utޖ%�i�Q�;~j��7�����i�[�u� �p�:�T�H|O��F�vuΏj!E�pkF���@�dٶԱd��k�҂�" Ԗ��jj��M�H�0�ov��	|��hF臵I!��?�0%�׿kҔ����N��ILm�~�`�R'ձ�Oz&�B,蒜�qEJ:BN4�k&�u�U�"sߦ���a 6�魨
6^n�L$ ^��� ���*�b�Fc���f,����b�N%�� )�(��~���A�Rd����`��ŧ�M�S�6�r��>��%3�j&i#Qt�y�d$S���|FhTH��v�������p�]^X���wΚy��T����
H�2����f�9 R��ӷLAM��Wv��h����U����H7�`�ex�G�L�m�3��@�Z4�yg��ݖNI0M�ml�\�nHn��۩��n�G�'�A����;�H昋�30L�'M��z�A+9��A��#�IBm��ڒ"���)5[�r�gI�jG�yߡ���(�v�ZR���* ��u��l��J*l����Dhio4�DI�ޙ'�b:����?���}�4P�3��L�ۍq��=�4��N��L&�7�&�D{��F3xܽ�ڌ��qQF����ܧU�#�Dlϧ��2����э�u� �JLmuߵ`rE��i�H��ͯk�E��� �:���b��8���oP�7��w�@���k�]w�J�<37��=s�10�m5�.�lt���6r��={Б���)�5�˚`�Y�o�j������o3FЭ��x�v��=�3�N[is����"KgcR�qeU���d�tp�L�W:�\CR`D�~���f-	u�q�L���2Hm�6���- 4�K�rfx�-x^u3|F(����U��2�56똖�ᄷԉ��HU�rI��ޏ��Iv4:�G�YV������8�Iao�?Tt$�3x#w�lM�-������v���T���t��4�r[�)Usf��O� �BƧ?�B�t���Q;ϒ8��%����J+��ߦ��ԄH�y�P����38&&�7��2�߼Q�U�{���kRݢbu�_٦����$�jh�L��I�9�;T�e�cYxͩ���'~晐m�{��q~�Bp��g�0�����Gy���ȑ�i����d�O]�J�&���ІUL�ڕr��L���?E.�:~�hvb8ޒw:f���).<P���Y�N�3�v'��f,����������PW5o�m��xD"sx��5(�{�B����e��kM!�o����c2i0�Ip19%׊D�ߛ��$"_9�K̖o�����]��jh6fO�M=2L�Yvۊ�#0��i��-%s�ۭX� ���`��a�M�oD�	0��F	��<)�҂`��v�K�!d���ӥF�,�՞�n��!�:ŉ���r�0��>i"H!�D��>��Vr�@� v:}��S�=yg��S�O�Z5��j��ۏO��m��N��&]��V57����bӽ�"��v�7�B/�Cj�Q"ӝ-ƶ�R�A�~���\�W�k�ZR�I_{��?-ۦ���}�|ɿ�@���ڔH��uo\Ji�c� Yy�;Mk$����qI8���ZT&-K���#&�Z�c��h��38��Q ���Pr������ jF��8i�M:ƼU��i��{d�2�A�f��������0,�q�H�阜���b�M���84q�@˘���g�;Z����H��6a�֐F;ck���H�k.gO�а��g��#����&���%���~ؠ�>����a0=����E�������3n�:�MW
�o��-3۽H����?�![I���y��YCL��;�K���sn=��[{��@aȜ�7���I�?kI�\H[2���V�W�Ҋ%�{��Ɣ�K'V��Ůg;�f±+x]{��+�˥�~h�_8��� &��x]����ԆW.���Yd��Q=���R�m��+�`��!�U��t6=8��0SK�ޱ��c>��Z�'�ѣ�=��(b�[��11�I
7?y��G!`����-"�o��M|�R����˥C�� �/�G4�u_kS�s1�_4���.um�*%k�Wm�!��I��ŢK�Db$G- A���PY�yc[G҄+�t�X;��)��a�؈�Q��b2.��Pq�����w�b[�� Z���9���HDT��lf}�
��� �PZ�<Ζ��ץ$a	�A�����&Y��i��4\Qm��fq9�FHg��(�'!�(� v�㯽dDo�B��378�~h�AȎ��"-�}W���j]ټ]��ʴ��ǭHE��Ϛ$����ύ��	���I=�q@��7���)�����rQ��:қ�u��C�v���	%V%{��#�L�ՒD�����D^"u���!$�Gj��Yě3�c��	`v��I$'��DL}�L=����[���k�{Q"��y�:��6���M'p�ן�I�P���<3tf΋x�,K��׹j	bh��� �գ����IW��
B.�-�X�45(YV�R	51��ņEU��� �8@��%��"��6$�MdK��h�F\�ZK i���:^4�b��[��p�ZA��P���.��eЁ��8�
��a����^ݖ�K$�L�;q�I�M�C1x�צ�!xf�2�MFp��
0P/��c�ďV~�(�'H�L�����[�]��:����PGKt��,��u��ߥ^W��R,D�W���lBBG�7�mP�
G��Co|�0,K������o���pL�/��W��q�_�ol%7O���bl̵p	��y� &��"�i�owքg.����p y�����k�ׂ�r�{t�����V��^6�ɿ��<Q�50LY���0��1}x��A��}��L��kރ���"�~�Sw�lr~�jP$�Ե���H�zƂ���pk��9���n�E0^#|	�"�Q�nS:�y��M��d�hn�G�D��%2�˗�)�g��Ԭ�:�[Ҥ�/�y�70�{fq�3b�&7���$�[�T�1�ˉ*)l�����MN��Ǜ�)��EǾgjC9lFT��2�Y�*(���=�Zg"`��t��v��2���K0�H����'�H`^#�Db��myV�V��-a��`�|[��N&��AN��o]�T����D���uF�������*ɗ@KX	݉WJ�js�~~~�eaA"0D�[*���)+@�v��eV����~V(�Zwm�?���,4sߖn����\�z��Wϣ��VP�r�N�.gq�*�֋Kq���j(	؃�޴���eT��,Ux��=o�	uPNE�޺�iO�����\u��y_��NBǏ�.I#a��9�ժ��џ-��:����C��A�D�S�҇ �?���<����|v�N-�A�[���(���� �[�ޮ%t��)p�4\�D�9#~�zU�c�>�F4U��u�ו9WtUf�	`L�D�PB�]���l�ni��r��?)�������V*����R)&NVs"5mt9��m����'^x�NR��v?y���m��2^�x�Cu����B$P��� gLf��ǽ$J퉽����Լp��	70�n�h��C�`U߄-y�_���:s.�T���[��m�=9[��Ğ(�X�ً�i�R�Fkq�{ԉQ��bbA���[�� �p���q��b��wP���lT�!�P�2]Hbh@`/��J$Y��zӢc��Aۣ��֑��/|6� ����]f�08/=)C(u�H	8�ҝ���hu鱽�?L|��bX�;�z�� �J'܉;"N�J�N�Q��zrh�;�.�!z)�PZ-V���|ҙCy�;h	(g7w�B�h�M�*�캥�h��F6Mrf� ~����#)��Zh%����]�n��"���zo?�i�f�m0�� ��� ) ! 1AQaq������ P�0����  ?Z Q��PG�r�����VӔx�TX�Ԩ��Pj��@�J��%����h�0�0�z�=7Q�N�/OE�q�h�x,+���!~�� ���&@W�.@��C~�f" �,��F!��WnlIT%Wh.>*���\ �Y[ .�L��7~� ��yc�*W��wS�����W�H^���Y}���l����	F
J�N�7���|����,${��v�G��շu4�3T� ��D�t@,��	�/\����'��	�0�e$$N6�ud�+�_�/b�`G��S��A�Ab�� (�%�煭�)E��qs� �jY�Р��89ZE[������'�們!14{���^�+���$O�D����&�*.>n�D�)��I�ͣ�֗v���gJ(����;L}ܳly��� �s*X���0@1d CxUx��,�� |!�ͻ�^�G��T�F$Ɗ�E	�RD&``r@*��a��˴���gE�	B-/�ltȠ��D���(��#g'L��+�C�|wB�T_,�|�\ 0��OA)�7�c�o� 2%���>:*"�@"�(R��u&�4��2��Mp���5ScMԓH��dPя�G��n���3�S�G�d�9���oM���y�WNβ:7���fj�K��5�o��R�4�� ���8ʗ�V�F�0x�[�tz{�y]��@7���4��H3���Bud�x��9����M^S�w��:���0��Zu-��HQA�e2�z�uE#@�H��S��q�aCϞ1�Mzh�vA9�˴�"���#^1ٵ4j�5������.��_��[�LX#4��E�ޔI�K:�и{�2�XNC��"����Y�P�t�7�	��94�j?�D�b
�Hq�B N0���=H'JO���&"�e4�Gv�"A��{3�T�^��:gRQ�J"k����X���'���h�G��v�ED�� ц�$r3G�v��"z#�zq��N{b �V��IU	��S��E��	<��̈>�����U"r��ݚ3p��ľ 'bJ�r?�"ES��1w˭5S���%Mm���}�k�3��K�j�)���P�Ab)��ݢ� �<.� �P�J���-,�J^/���%@(O\0�T\mB0��"P}� �a�6��&00��"�W��o�uːD�%^)�6$r���{'� �x�f�"�09���Z�����wH �<�pf�A��y>�N�M��$%*IU EB6��I��AN8+�Q�N��N�G�$ �MU_�6�4�H3�~k�Ej���<�q vR���6ꮈ��6 B,��M9��G@�Vr2?�u�oW1�W/ɼnt>�
�>�@`N�mF���	ձ�H��q'�/@(7�V�I�Ș���B!x����H2��"�p�qP��G�8Bi������È�a�բ��LGGw�b�)1����!ClC��=���hD�;�i��O� ���UY�8^������������EG>��l���+���'�;�5��\�+����u�7� �g��Ҕ��� ��b�w�d8�j������9��W>a�S�b��-����%�ߑ2����9d �"���t�܈�MT��m��ʽ�U�I1 5U��IM���z�J	����9) ?l�aX.�é G+�#j�)�I�E�e�������r�F���+��.�
��5�A��]nP�F��R������g��^����ZF�8�I��B�o6P<���/�\�7�S9���u6ނ�>�����k�)X�$F��-���X8��)��*�͖Ƿ"�"��� I:~:U��Z5:j*F�@�!��+q����lx!:�,�	�S�1@���2��<A�@D��%��R�J�/��ךD�b�DR��I�&��:W!��5@���T�	�v��#F �9�Gnʲ@�IE��=5�6r��Φ8hxغ�MDp'r����p���5`���F��D%���(�q�|FT/�XxmR�SW���� -�i4�,��tŇ'�'# (<�$�E�8�J�JT���\��0�m�A(���*�����E��5��r��H &bl��p}'���J��Ҩ���ʫ�!�Ri
�5u�!D/,�%
 $�ío��_\0�<~��=n��`�ï�Y;�^�rH�+�t~ڪQL"���xt�ocd�]�>��x�@#) q-}fx��H�����^!�M*'��*eV��B��}�<�w�-PC��#�\�$U'����G➽ռHi��d��N���.��0�����)ݵ�Qoh���7Rj�L��8���4��j�^��H=|\�J�Q# �*���f���Z�h����"�bs����E<�৔!UjE V3����I#��<Abe$w��jW\��*V)	A,�X�6����r�����	��"�(�=q�&U��5Pf�g�ax�"��=��m��3�-<����<:��iW9;�y@ �r?5�C+ v��4(6J�@���	�WPg'0���b�(�D�JETd���g�WP#@�^���ڕ�	\�);������_t4�	�Gt�Dz��P��"�Iy-�8�,2�����
6���f�4%R�F=�C�;�s$!T� R�u��)���7�j(�)���� �Z Y�E)T�JX�/t@���QjG`Qr�>|P�C��R1/B�Ye�$��[�:FBq}�j$��	�ܓ�Մ@�b-��֢���p��f	y� �a�����X�Z�?|� �� \5$�7���_Z~�<1�	>���"r����2�˝-0X�[�=�������>����f�L�D I���`ŗ�d��q��XB=�U`層�~��Z88�OEd����+}�f���r��ݴ��TE$~¶�Yd����Cr_�ԩ��[�Hiß�fjVc��sC\��9:�O;AF�D��R�h-(Zq�}�P�)�4�=��Ș�ˢr�$#��u�#]iR',�x\�#�&�H(����-6|*���ގ\j�	Y�SC�+��I�Ȑ�L�5!]�R���A1����0N����H^qQ�9�� y���Պ�����qCp�=�����@�m�~ �B\��@� �=DXu��E���n\H!&�sm���W�A�k$��B�>t�-��ڡ� dF�A�2�9m�q�C����/�"mt%���v9�3�q'��X���"���CM���	;�F |
j�h�# Ҍ+��	=�,u'#t�*[X��8vt���=� ;@F}�O��W�-� ��5���8y�{�\IƓ`�ڜ�h�w�Vҏ��,��t�A	�|���*�d�q�w_\I�W��mr!j�C{:��t`$/<��:���3ŋ�IF�jؔI��Lh3T�e���A��u���iD�F| ��ӫ0p<��Pe�W�X5�vMw�/�'	ȹ%�
�&zG઺ݓo�����8��G��3�v����jQ� P���4q�����M�������aZH��5�@�p|�oD���KKPQ��f���f�'4�����U��x{��,��hT�K�4�A�R��-}� �mU��#��ߓ�����_Oop#<{�ȯ�Թ��զ;m�ᑍWXp�i�"���J
�@ 酪ǿ��^��(@p�:H�
���Z���w]?<��/4f�\}9�q[�é�n��|2���
$��
H �h�UK��M�J<	k�0��;wGvq��^��m���ц�`t@�YO�i8��nn�=����J�a�x��"����:��/��'ƊЭڌ� '��T4-�e�
��ޱ2�u�<�)��t�vc�*�)$n[FJZ�#F�������>p�1�f0�D,ߊyn�6�����3x�:/���ʔ�&��Ry�v5vXtBq���.�����Mx�7&8z���Jl@�*��Oi�� �
�����2'<M2�%��d�
�G��|-�Ϊ�3.���{ vԼ���+��ǃ#*�a0�lk�v:�������[��d�;؉�lXr85���h5�а�S�t	��[6�8JE28����2���������E&���*�e1��տD� �)^(��� �8:�M�Tӈr"nHȅ{�Q�5�*�͗r�]��P�}�w��<�;R�ir���AT�e<ʏ5�o�%!i=�:E7ޛ�HB��n��= ݜd[�vQ���2T�Un � JH˃��J�F��ئ�	Ҿ<C*��A�=A��\����gpz~r�ˠ
�:���+.�}�N'6����\�u�1:�*��t�Sx��[o�m�U���S�1�p�hPQV豰��,�(
����ȅ�Ս;%��d��.���8����;��fG\��	�s��ˍ����@��!��D��>��݂�U����mH�>¦;M�]=�\@/�,�b�!�H���sU%E�����m�
ag0�=s���J:ď�X�4�zY�.m�ee1�}zd"I�($B�Z�S)Z�t�2��h�(��m�;ǅ��n�pu��q
H y�n�N��s{��?L��Bb�Пꓴ�?9X���e̾f]%�
�1��>nN��ؠ��B��p��A��h�\?��1�F��X�L#�ʣ�-+�(�LÄ�+�SE&����m�Vعȥz�}_(��b�Y2B*�Σ�T'����[�5�57��D�JD�@_Gb��qiRcӝSڨ� |K��+\�k�a�����f�Xj}�����@K�pK����i��
�>,+I�+vƌY ���:���*R&ڂo�pύA�5E�`�:;�*���:�ᇄ�0`D�ʐ����/�m��xߘ�|�D��˜z���ڴ�9䔎�C]:L���;���ىu$p����@����H�熭� ���b��pg�ylu����58�
�n�jR,��(@.�g��X�W���~&���wa�<���k6� ;`ŀ'��C8U88��ܮ�b�D�{e6�Z��3zB�C�@T���0l �CZb	�8r�)�z�I��6��$9��v������&�S�'y��8�T4D:�{��:B�ڨH���L$'m�J��Q�;�Ğ����X)mT
���
G���|�Rx��;!�-��L	R� 
�S]��0��8���S$=l3*@�A;�48�������z�{��O����a�d�\����@K��1ҟ��nX@sfPMg (��q�ʾo�=�\�@fP��ʰ�g��~4SѮqJ�Ż��3����b�6�kJ%�U��2ڔ/4p�#�]"#�@�B�7	� �15Ќ����=n�P�_�1�����R�!;?�8L�|��M�x�gY�90egBT�g �������LF�f��ͭ�Z��`V,��&IF��M��}����7�����]E��i�$������yl���<!� ��*��(rsw�:����d�"��V!�ϻ�V&��9a�Ƅ^U�g�6�0�ձ���F1��"G�+�(]R�8�ʫ4��h6�+�����u� �&�Y�NOVV)���J��T�g .=UY����*�@�K���7Q�K�7�������j9
�C;;qk�/��1|
P�̃ �?���Hi�p~_�t_��)6Ur2q:'��T�5w�b*	 EC"�)GB����������g�g3��(�v�,7Z���n)�b���,���H�8P�O�l$(]k�<�b�
� �+�>�_v��R�� �b�����AT��<���S�ƞ5���ժ}<aI��I��U
N�V)T��� �rh����yK -"�M��)�r�5�J�&�BhDG
�h|BA� � FU?�<!�I`�hã˺J��W�y�Y��.��X��[�z"\:�H'gz�OG��+�z�n�������6�$�C�غb� �sW�>7ؿzY���
X��4�	�f��9f�
��P�eP��TZ<� �
�Bu�� ��IS�:0��ew89���7�y|Q����艈7�͔V=��6<d{OZ��G܁�9V�pxłOP��G��TP���1�%:B�П'W�$"�̵�����8H`��UK$��f0Q��LR�,�:j!R0)�{�TWϑ��ؒ\Gp���vb�� �`!�f�w6V���[�1�Q�UL ��u4�Ci����Q*˛I��wxK!Y5w(�����`h��E�æZ�r��Fm�&��/I`&��w�V0�+�b3«H�4o���wF�O��˓��|A� ������4�
�x>�<��X}��c�و�н�p�?n���#ܵmB⃦�l����jo���Nȝ�9n��>�_�@�:3�^^�$.�PS{�F ؕ�ݘxn�\O2�D6�xT��oy���V��y��!������W��WS`�� &�����R�y����MWp]0���
C�� g�vU�J0�Jщ0��!��@pϖ.E� ��o�]}��W��aZ�(�Ȣj:���$��ETH�%��`r���P	4U�i�G5M�L*8R΃B�<hf���K
):pמ� �&��&$BJPմ���@T�3&���s��B����P��kQ~M}mW�ڇ;�O���8�d" �BN���_
�k�h��^]T$(���\1Y/]LK��	4� Gs2V��R"�Aa�ҥ�n@E(ƈ�Ě�t�օ��-�N��3�"N6 �����r�]���� ��*8M�� ��!���l)�G2��^R*w��lJ>�r!����E��.��r�S~�(��,Kg��&�iM�䛛�k��?�f~��܌��u��Bu���T=�I�A�P�Bu*\�K���%I�����|/s͉�)�A�2* $���	J(���I�M=\^�	� _P���t����|�f���"0H�H�O����6�{�?�,���=F�������灂ទ-��U�Y˻�D ���):ЦyeH�[�$�އ�$e;��+-�qR���ɦ)!%�d	�< k7�)��7�7��J-�������a��qA�0tL<�Z:A����2�gd��D���IJ����L��'�W� �0P�
T��4���FS_���|ES����O%���!���(�+
�@ ��cM��ԁB� ӗ*h&j�����3��FP,R
���PBĒ#�@UDQ�SО��-v`��|�����	�G��"�F��镃� �hMUw�>P�&py�آŵrJ��9�)�-O�*���m��8P'E������8"r@y+wrؑ��TF��6Ð�K崈�]X�\  ��t�%Z�Ս�0[���o�5�ƣymCpH��� ��QP�&u��K[1Ku!���{�m����C��0���AT(�
�X��E�8a���k� �I�.�?��
[g��iu�z2:��d��m!��f����x*���V/�H�<.����o`!��IJ �.U�RG�K��e�"m�~xbD�-��G'�G1��-^^X��3�pb���C��P��^_��JLmG�^�I��F�W �y��"N��_U�H\eC&��H�#�0gL�)g�1��h��W��,�B�J�	I?�W��S�xo+ �:�ԧ���$D8o�|g�s�n݃g�9� ��9�p��=P���;u.���gdd�ˠ�:�xcDѻ��U�Y]1�lڔ�~O�b$�"�K�Ӄ�s@��1��<d�Q�	���9L�ŕ�N�@�p&��R���� u4s������9����]s9��@�.�yur՝�,W���	����)^D蔉�!H���UR�Ȍ��@+�H�I���u�p��Q�&;䟺�UB4���~+-0�P�U��ͣ���U%U����0�R�;����My:�8��
6�) r�F�*[�H�"%E%��ZM��)N�T�L��O��N[qZIraj �1a�G�M@
%��P�� C�$��)�l���9���PIhC���.ZLB,�� 9~z�E<*J� �&}8<�;Ǎ*-Q��{�w8�`�6 LM�""����ߥh�[w��,����`M�E�g�hEhԐi���IGH�
�J�S�jJ..�8�/���7��yٝ=SG��e|�n7s��d�n%C�D ��:f��`���̭c�������ꙫ>Q�_��PQ9RPK��`rH	�!�"8��+s6hH�T�tf"B�(Z�H�b�ir�$�o�Z	?
�W���NIxyq����XDu�R���@��Z�|�NOY�>�%�g������{,J<���hh2�p.���M��4�o*KH��'<��SH'l:(��[�e���HT�Z��L@H�z��Td+Z�_�|-��L��Z��%���{���T"1�"�T4   ��[+B0H4FC�^`i����<Ĉ�e4xE
���mT���ZS��hP���1T�E�'�� �L�^�uR�XS�hj���bx`Ak_�j>V�}� 8PЖ�R�Q�"N�GCk�$b�A�š�>)"�Yúw�<P��p(�^�#�X��P�AJ�<�� Ǣ?�o�� ;ev%j�(��'�BeTb/*���Z���o��q��h<�	�E�hR�T��X��N,!�ձ*$s�\A���9H�*,HՓG��Oɉ%��~@4�����QQK�� j_��c�(�l_������?�`>����J�{�f|��pMZ<<���8iG�OB�����t��H_gϛ�/���Z�n�ǱE��n�}/%��;RP W+�A�)�SҺA���y�ƿ�"��Pɨ�x�~��gۗ,Ԝ@C��H3���|���T�]i���E�-C�L&&_QcG�4�$b�j~� ǚ� � ��77�&��@ ��������y1�4x��MS{�������S��F��1Z�1��c�9���
izq�ƱS���r&̸ke���F~>���Q�wݞ�5<���"6�e��%�(!�"�áI��QgZ��/'�Up�7��Q���T�F;^�\f�O�[4R��2Az��gL�+PCs��qMo����ʜ@:-���~�dD��/�}ׁ. 5#��|��|8r�G�J����c�|i �o�u����'��	�#矟À
�\Q�i�ڿn�"�}���x��bЁT� ��e-(<P��6���jPj�� ��u������S�ߜ��0�RSQ�O�D�
K��@��f/��.֕>=�1���f��IA�j2E4E8�N*&�D�H8/�,���`�
���*�.�W_3�UQ%9_%����v/k[���%P���廞�i3�+|�?�*~�!(��lʁ�V��[>���랓�K��O���� R e/z �E���:��$<��iP�o A��������j��,W�FL� �ޤmP"�4T��]����D!T��� �;� m_V����O�r�<����Oއ�?
 6�*$C���=��#�M�-�3��!�!@u���Ӓ���(�{�"�l�B+�&c�=�%�;��S	3�_Zr��OSF�߻���L�A&I4�+��f�$���R'�O���k1�:�M�8Li	U'�z~zB��j��� ���u��	t&4`�.�!��,l ���о�R��rViє���^7Y�@e<��T*������ �ȸ�~9A*s�gACT�f�W�A9�x�#�� ''��H�8U�'H�:-��Ti���ܡBa���q���c�LeO~�Y��� p� ��OAj *F�h7�ƨ�Nzh=���Hϲ~�8��zz��8Y_��¾:������LNS���iWV�e�I��s�X����H����P���@0� }3�J4��� 5����OBx��������$�~rP~5�t�7� �I���Zo�bno�n�j����Fo�5�(�ш�����L�u�5�⭤�n������-]ۈE�,N���(��*�e`���T(��y`aO����Q�	��9�o����
~�vɋU�e)�5�V�!�(_�Q)��V^FMZRЇ�|�����g«  ���������x<Ed�U���e������I�F� �X����m}��`��P�-���V{�
�Z�B_7�~�+��
��@?�H*�us�#R~��&KH�� S��XRcS�R}�)E
�/�j0:��S�W� �D�x����*O��۳�<��!������3ݛ8��9n"�M�X�ЬYI�B�ӑ,�]6�r�Ò6:(2S��T�P/�Xu��b̉\����M	�����l���v��3�}�#�>9%�@HGVJ	f�&Pa���t�u���� �?�6��I�
��Qs��eU��� �_(#����6T+#F���,����$�����lSf���\9X B"	}C-P}�u�Q@���L_����yd1���N�� /Jל`	�ؽA�G[��ғ�;������P����ߪ����1%T��� �� �\��C?������	� ���n{� �J�LV,3DO����`��p~D�|&�1|a����C� �lP6I	�4� �̡5��B�����p������ ����&�"9O��|� ��� ���ס']!>,�X�� �/�����Avw�&�v�Y���b�%&yVN��bb�=�Ņ��47�y�QR�s��@�dlܱ�D �5�M@�;���?�(i�P���I���Jb�v�eiQƴT<(����ã$S��	R_>g�|#������0��)�E���+�����C���sn-6$7��Q���������!iBU�_�� ��Ȇ 8�U���T��P�pv���/�p>� ��?T�I�(�j�N��=�=�xt��9�i����3?�jIך��;�}��`t�s�dW��	�����S��ŵf�`�\�h��fbC�>.0+g���>��h���bYH��F��)#���� g�돆�vAi�wP����1��[��=�0�dU���¯�pP|-��&k -1R���P���X��>�I�"��Z�ѐ��	�����'�o��Җ�AQ� ��y-���&��mÕ�
��� �/�6Nx�t�j�7`���5��{P�ɔ[���1qBo���8�[��BJr��E�=F�XvM���&����x�!�j ���.�1R�t���b�W�|����'��� �堉J�~��y0��dc����aJ� ���LY�(hW���d5��h9����T/�c�W'�;�U��2�� 3�����g�-u�(DjЮ����^���?��c���^���� Q$y,�G�˝V��
��$��i�@�T��� �@An���Z� \� O��;������!.�Ť��y��T�l�H�Q�$r&�ik�zN$��)�E#pbtH@�]�	����JZ(�A��x� |��-z��)�W�������PM'K����l����[���`��ZO��V`&�R����_*������z3��� ����� T~���?�y2@�c��"<D 0����[�����B�sĴD�.9����v�(��c=���g���aAf!�P��������D,ؓ�U8�&�+ ���\�^�y��d⵹�-i���-OC�B;�����:�a�:S?fXS�M�La�0�P�p����;# ��؃ h�<,���t���$A�  &q	E�)R+�c[��BQ�++�_�*蓥0 �j$坸5�jڠ�Q�2�3�!���CD��0�Ȑ-l�槨�I��bdj�;�}�c�OM��R�b�D�ߡ���+�A�Q�)-J�����L�Q��������U^@�0���မ�/g,�2A�p~r�b��I6��K���a�7��֢x���_�t��#ӏ���f���6�[b�6�\��6���~I�&�B"���r	!e�~˵����T�-y��tq��J���8�y����Jg�q!�d��*��i'f����O��ԛT:2`�t�,m�^��6P�'�'��}�1NR�3����^[�l��\����|k���?�#Ψ�'���;��^�J����3�a�c���n��? �w�12�F9��\$������I�w-�����	�u�<~��X�?��������x�9�$�#k�/�d`�T��X��q�$�Z1\Wd����ɘ�I��~��=�/�iOD���2ҥ��&��a8�
��b�U�Ha�M����!Ml��Dd+�����$�U�X��~��ɦ�!����_��A�&���d"�r	GH�RU(�W�66���ƫ����F�`�77K|*"�}�1�}+���4wCX�!�ë�I�ۛ�N??K��]��@�~��/������T��V��0.؏9*����?����}]�{#ҷTu�C&ج����<���+��t�����T�Og��40I�z
9�Y�RñUU��y�t�s�����?�ҫK�hA��\�^^�^,-\�ڱ�lk� -@W�q�T��������8zY�Tp�Y �c ��k�J%���	����;�N	�2%lmr�Ҥ��vc�����'���4�LZ�=Õ���V��p��
����q?��;wB�?������x&�1?Fb�,(H����WșI���5%�OX���ʈ�(�qD�S��K��@ƃ�.���e|��{Pu����[.�f)�ߗ=J��6;�0��G:j'�%����U�������K�$Iܢ b�}^i"��t�d�4x|�eEQZM�]��������?=���U�h&�ޛ{���D'-�����o������s��Bj��|�O�Ak��9�L7�`�P�V�3{}��s\���	�q�mU���?��ᦴ3������C�&��c���g��"�J���r*R��ʟԇ<kף� ze�D��!^� K�j����8O��h�3�ڻ<B:64d$w �J 
?Bl��%����:S�g@��'q��S�W��D�X�h���	[�Y6uɮF=a����E'#�m�Z+�n���.Z��%�4Eb黡t�����^�p&L�$��O�����tbM����g㨓�F�*A�U��"��m���}	xH�',{��!��t}���2|4�`��:b�

��2��+bF�[O���y��7�Z��/�
A����[�ПU���ۙ�wm�tE7�ޏ�h(k��δ��lrN�|x�S���H���u`�������$���p��s��*�xi�'U��p�8[�x˱N�YL|�;���b)���$wh̔�rP�#�� ���0"�	l �U�93�1�\y�? ��3n�}T�Q:YVIi2����R~&*җ�ϺoQx䋦�y�3�~e�?�6���V]"a�<�\�U����X�XX��<>"2��!�)L2U|3a~Ѣ,�W�l���fi�N_U-�a29�*�����B���A��@�8Rz��ovES�7�d�(Q3�j��1���E�ʻ�����c�����|*���%7K,�n')���aE{�ǫ�쁶�;�w�>b����L�x�@L�m:�Vq0�$��*R>�g!����pEb���w���|T@��.��L��~7Ui���3Ǹp�_ܷ�)�������z�`���QT�aj��_&�2ަN���'G.56*�e�/�ɕ�� �[M��#Ǡ%��(.ޕ�I@K��¨�'�JS����(����b�[��*߶c���V��44n!-i�gy�q��@Y/�Zuܤ��n5��O�\�m�.��1�X5�U/�LL���~=o-��P�~��c�EN�ԍ�w���Ó�hfO�u��޸�g�o��5�T%k��R:��}�UW�6�>~^�&���j�Tu������X��Q�������H]g~�b%�ѯV���2����fV�uW�)�B�_ׇn?�s-��\����W��C��b��_�EW�(Egk*�������CAEy�##�*�l�*.E�W�<f5��WOW2�-?}�.z'��G��_ͮH�<�tuŽK���Ӗ����
��"?g�uU��(>���N���PTM+�<m�k�i䨛�j} z�B��p�u��^=��\x\0�{A�%����#���wx�
�.	��U��uz��������WA���Pq�����s����Pg��a0}���~r� �&���3E��X���$����f��n��ƴ��PE��L�G�@e�]'n,l�)��VD��B���@bf��A���6��%xy�-���wP��yЇ*� ���aod�����ͅ?�f����E<`��ᕮL�K:�Rƍ�W��1�,&�n��>����Q}<8��04�������x�-y�_�"��ׅDϩ-Ô�L	H�%�z_}���֢��lf�Tî�G(Rdz��4�������:Te:�+qVEJ�����F$�s��s�\Zt;��q�3sO�_-ۥb@9�W�#��+���mk%ZG�[ԘQ�P���Ǌ\�ruK�vR��cs>�W[�Z�.7LD��XV��C�M�&*�����~�U�����*��ݍ4�O�u�Ԋ�4���BWx�ja�[v M�������Q6p�_��Oh���|U��������x�6Wj�~eܬ�Sr0����ֲ&�B��F+�n1#.�/G�b��鴭���sK���(*�+�6u���kyl|���H�^�F���Ɣ�\�e�n_QϥdFa,4���͏Cn�&Y�_6`�>3ف}��vV2�=8D᥺S)'��[m����@*�'	�~-���FQX�dޗ�S�?�(\u��hm���3�Pj.�O.Q�p-nR�~I�f��\��D��2��f�H���g�=��{{�t���Q���F��%���H��\�d���g6uT�SkYp����X�J�o&D��U��:�s��X�H�W@�K�sCb��m��Ҟ� d��}A�f?r�r��?`H?+�����hR+���6"w�?�C/D�������B��y�6�ۇ�}FG��!rL�j	9�'��ex��T����>���[�� ���}'��Åe�<!����	,��K�ꩤ��L��w1�A�ƾ�*�g�E�^�R���#W���K��m����En�
��~��!"C�%?:��W�z���SO�tZ�̣�kv��΋+~��]:p7*�ngr-�PG=Yyo&�>,?���L��Uq�� (��w��G�Ӗ��ʕ���<<?JB�!���Y�짟����3{�O �T�nO��j�P��1������h5R�gu��]�	*;�N>P����_uvx^se��[�p����j��<k���\���>��dμ�ˌSb��E?J��8��y&�����ǴH�s���K'�9kVׂ6�c���R��+{�_Q��A�n��*�/��l-nć�$̤���Q�F���1,w
P4Ԏϵ��r�
�$#;u9��t�rsC��2 K	��7�l��{���Ոf�����Qd�=�W�N���4��H�~����U�r�λ騦0�5�35��r���xC��G~�,�"��fOڨ>q�4�Ąh.�a��*��Eoǭ�����$ҝ3{�p6��ٍ�I9T��Uy�~̤|��˗���Oh�q�&#���KM����w�Ưl�n=ϊg^
P�H��ĭ]̷:!0�{��Q����6ORPA��D>�}�m��~ȷ�Ǖ��~�E?Z�v��}NSI�(�"i�?�@%���P���W1��Q��5Zҵsu=�dC��x��l-��Xӫ]�N1�e�d��Mmc�R�r�ء����}{�PH�j� �Z�lh�� �p�(d��T�Ʊz��|�p4>Ȥ?�xe�A�sd�\پg�tb�v��g{2[4���3���.@�h���_877�`hL�΂1^���@���Tϴ ����A`�%�������"���j�>�r7)���0pV=u�4�����k��M2��b��:S�p(��ȩ7u�`:��#�6�
�c|~ 8��=N\/ON/�}�Ae�q��]~�h��/ l�K.�OX��٫�-�l�0���WHf~��n���Mt�^yhS�'�c�r�m΂N)���~iv�����t�"��&�v�z>;��K4�����{O��y�00	����4�K��@�q�)�� >|{$Â�':����.rLt�w�ٟ5?'��<Q�H(/������\�7J����(�6�����9�~_���! Hu8Z��?l�r���8��g����{�-I�|Ş��:�%�*V�'1hb1*_�7���͸ 0H��D�vo�|�$zw��Y�#]�"yN�?�W9J2qߏ0�����5NHC*W$~��:�ޝ���Wr�^Z	��:�R�vq}�k��>S~	�7�a~u��(I
����mC��;'�hhEҪǮӪ�D��n��fy+"F���XϫN^R�!��_�>t,����U�S�O��O�[�L8,Q>��y��G$>?���x%`��`ZY�oۭ��̩#' �MIE��1ҍ
UI�?GtLj�a�2<-��jv�-�,�������$s3i>��zԁ8�����$z�����mdI�V��UI�4�_�:�0C��pMiN��i��n�Ԙ.�x���ix��}�q�c�4�;�'FH���Δ:v1��q�F�u
� �%�96JM�J1��~���!ʧ<�X��򘺀�ɴ��P=�J��.Ȅ7��l���S�q�x���YN8`���e���Ѵ� tэ�NF��m�͘�t��0A�ٮZ��f�ZC�)��E��Wx@A�/�Y����g��Ӂ���]�|��E=ٗ��,�kg����<Uu�V�{,�N�xC���wuENAW ���\m��3Ï�		�Nv���D���؄D[B�'/j/���,k�#6ȶs�� ���*�g��>��4��F�d6�n��#2��ٳ�r/�����}�IJ�.��̷�i��K�k��$(���Po)�����L����{^Ȃf_��>����5؜�
�Z�DL�7���t���[ w�ؓe�Ο���?�J���O�q����pG�{���aD_?[��9��#��pj��8"��0��m*�ص�>S2&c)i����i� ��n�x��ګ�������ϸK;�x G�mI鵔:���7�<G����lS�l��ų�;� <}��!��l1�əA�wg��|p�/0���?!��DV<]������b@��ݧ+uDk5^�)��b�q�T=�CG�`n(���j���o�/-�bu���\�W\uuD��I˅��� ��>[����=iz���:�'m�?s�J�p��Z����@LU�\���l����e���������'�/Ί���W� �Q�����5OS�.S)�=~�k7�<��I��W��)?������}�(��т�)S�L�=��p@_�Ȣ�DF �O,�'�q3�E�(tD�����С���R��R�q�|��NWFh�vF�������W������a4�ʃ��ePA(u v��l��\s�e��tTw���kT����C��-���Y�Ǝ������8�����`B��չL-Xg!> �U�x����F�>���Ry�M���v��N�{�]p�wYٝh��򚖮�UQ$m�B�<�N�Df�HbX̺W�Д*�Uv쓤m�u�F��FC:G+d�7g��_���%�ʬ����N�i`>�O6y&��|���Xk�#VVq9�~q��|���\�a �W�^���������!��t��$��iH)�~-��wc��"1n[��wGC0|l������� ,�T����}B��}����\��a���ϩ�2�d�CԱ��	W���-�������� �5�׋uQ�A:��u9`���V� -%�����|�|��/^�A�j��� g�,q�Z�R�������)��H�>��%��w\�����XL"���I5S��ɨ̼�u���B-0��cV�	�[z�\_���_�_J��Vڹ;�+;�8k).����h�X�X��ȅ�(b.X�K}�6�������b6Z0�2�t��W� �!���7��#.���Q�IHGe)[(�`�{���3a�~G����Q���(�_4}��IB�2Y6Ku�e�Eir/<���HנX跞bʱ���.��5��$�u��ߍt���SiG���A�41� �~�C�	���f�*��,�aU�W_w�XW�~pgKx~B�X
l��d�+���b{��|z�VyM
K���a%Y-�4��E�׬R�u\�M*|:NB�l�9�4M��{c��7h���7x�K�	W�k@
�?�c�8���yX\��̧٤;��g��G����8\ōd�hF2_6���-�V��_7K;j{%:�1��a�z�������Ǵ�/`C8�?�B�p h�e��C��r)hc�ɕ��+|�x�N�F7�5u�;[����?�Yr�o�	��D؁�� ����q���ŕ�Y��@�$pB�J*�:n��g�D��[� +v�u��d�gra!VS�t��dd��l;8O�p����N�8��>�k�C�z�Y�F��̙�0dꌓE���d��y��*��-c���n
)9�US��MK�w|�)� g=��ݟ��CN��|I(ŒhkM�Z�d@���#��#�"�:麴%&�@v�U�k1Hwv��!��9�r�L2HNB�ן�e@I�5b�emk=Yv��K�+��|��O�/	���WT��$�xi�NG(�ݺ��heA3T��L�;j�~�v��w�l1EӪ�FE�\F��LG@GL��U)N~�[��N�@2�Į�&�wGOV���ŗi�]��ܽ
]'9ͥr����p��{��9�Ͱ\��oCq;�H��y�˞g%�H�7�GlԎp���U�����^"#̉�"�܁�g�V�5ۍ�&��cTW���53?R?���%	�.uJֵW�Z��a��ZLM΢B��E�,��8#��V����ԭ�J�p5�I�A5ڪX�Ok l1Ǡ]2S�U�M�o��>�w$/�x�8WyI<� Uf�,9�u��l�MI��]?�{���q:|Z�H=N�wu��r�B3�-��Rg��������V�cN&���`Q�"�7A� ��F}���x(}��<p2�x�� 5髖��D�g���s41W&�t�ܥN?��Q�E����c��)g�^��e�|;���[��2ʃ���][��!�JAHo��U���Dݼ�T9�����Qz9~�H�Ё)I��ӡv����kW4U@������J��w"�piS�@��}���*>O������kwb8�O�a���_�i��`3�V��]�b�X���R�u[hD��.�%z8�U\���21�n����ܶ�ܰg��4iuAx~.w?\��#�	�+�+��d��1Z�C���N�
�JU~�͵�9�r���b ��h��8�Y��i�3��pp5��S��w���J	8�鋱Va���*�2e���Z��� W�/���h;�^WIŔ'th��v��@'
2�����B�PW�.���q��}�	X}�c�%r����w��]'s㭹����rj�r��d4F���7�R���'��w"��]�V�i���p��]sn�g���A����-ޤ熘R�/�n�@b��@^��A1���ș�W�Rҥr��{߆E��}�{��YZ�F�+� �O��μ�I� �1�Z���<[��\u�9�ߐxb��ß� Ӵ�w��!r��5� q�f"&�+�xS厺�X����kLi�ܭ�
�� F]牢i�.�wB�ز������,�? ��g9��"�$�%t�)��uaZLbѣc��9���GNnAͅg6��i���=o��`����c0��|`XA�m�g���R��~[��Y��6�}�)��oӽ/�c����hf�	���m��ü;�t1w��]h�ܷ ]?d�H<�O�0����SB�5�ȣ�Y�F|Q�ِڿ9d%�I��\f���h&�x$����H�K�K���S���\�'I�d��������֌��u`E�(�r��t1ܚ·���p$�.�w����!���;�*���<�SQ-c�/�nޕ�[*����R�=�������R]�H�6�b��.!;n���ɴ�a��tU�<8Y��Tk�������u+���gLD-��@7G�V�..�S�W�L�a�-h،b	��<���sTEj�
�V����a��L�I��	d%���NT�R�%�.��B�Mt ��V�&x�O���EP.�e�fH/4c�� 	Z���0QMh���͏l9r.Y��$�z��E�s��D&)��r����~pO�Vd���p]c��k'�sj��7hI�c�1��gh.*"�#Լ����,�����ԧ��~mm���/��Or��it���E���@����cG�
��o-Aҽ�В��kc������Hٮ*�q_���}R�&9š=F
tG���/�h���-�E��
-|}>�U�����lsVw���l�:WV�!Y���ce��58����{z�M���9�L��W�q5��~%�j�^�C%��̉PS	~9����g)�=��S��-�͢s��I	"�pv��iL���@�u��h��?9*��F�,Y���--�B�}�9��=e~�Cp�x���c_������iC�^�dуGd�����`�y*+� I�W�^"���{y�5+�Py3���~L��3N��"E�\�����x���su�]�Y�Y�����e䣁�S\���iA�/N����/ᬄ�5_>SUr��4�7WM~i���{L[;���t�����=�#��D⅛��W�g�6�g��c��?��h�P=��9HF�g�r�C'�-����?�0�Čl@_��T�=���{��j7�ug�?����~�q[#�׺�`-�0��͉�7B�g1�r��������sC>:)O��`����*�}4fBP��Q���n�nn~��d�� Ea0p�?,%C�A��|OtwY(�dPQ��6��_���׼a%µ��qK� <������q��%q&���ڝ�����C�)MJ�Ԛ.�/9c�2��Jla>�i�s(���6ml��22�j���x���G���/��8�ڲ�K��F�!���H�}���14����~{�?@ѬM�fy�����`I ?{��
B��nk��+�̆5��N-/�����1j\}+����ogՓ� ��ds�� �~N�^n�pF�o(?f��r��W���B�`��R��NTN2oPA�k�W9x��.�Ѳ=�m"�q�c;J[����n�ww[�Ol�&�椨����@(���m��)��ܑ�,��Df/}ͤ����x73ts0�C#�u�d���ܲ��z��A�ŋƕ�D���o|��E,��u��(Ab�$Ot!�h+x��N�Qp�>o?���s�U��Nu� ���(�40|(C��`�~oMA��&d�	#�2'N�X�B�$o��N;<Ps@�J+>y�5AW�����Xƕ$���~��4�-6����'�d�m��kS�E�{����~��j���S_�U���e�Wu�>�F}��x�Vˍ��d	lO���l[L��|U��=��X�)螓��P��n*�2�Y����er;[�%����|\}F4~��Y}������Rh?oBD1\:u>1�U�,'���D��	ef ��geJ���{�z�\��Ѯ�)�U�;D�J�����o.��2�~�����s%�6� ə�H$�&,�Mʱ">���Ze��ͻv��r���
?I+׮[�o�
@���S�Z&��V�;;�<�A[��g�ha���"�3��!�S�8U�Rt��FNAw�0�7��wÅޠz&�-O�/#��q���i�q����c9������eX�䈻:������$J�f��#��j$H��$��̚��\�R���È�q5�����L�rg�L���Y��q��H�b8��F�x�Qv7����a���nȌ�zZѪ�d�粌�EDJX��?@b1R�Hȹ�
F&-q9/�q�&K�����2
�4G .]o���`ߠ,�J����K	7�UX��=����_u�[�k��5��P�5�1�(�&Ν�Tݡw
r�5�AAq�B�8�_��Pmʪk߬��r��u��­DZfd���4�ى�`�l��1
��dR6rI��63�{���}��Յ�&��r�9/�wU�=�Jqd��\��-`.�����F�X˵��V��Rr�K��uz.��r0�/�)�\r������Sl�C�wZ�K2Ѩ��өBk����Ih9�mN�U�i��p��5M\���<�z��8���?Öcb�:�;ݽ��y�]�(�����E?�
�G�����ۢ�ܨ-g�q��	V� 2L9� 1R2�f'H�@���e]9	al�jՇo5���+���X6�7��".y
bY���o��G��)żq���aoC���藩:ָ�xQ�k��q2n{n�S�^Ec��1����D^7���Gi<�;+�,Qb1��Y��C�Jz����@M!d0���KM>��+�r�@�)	Ow��E�Ŧȩ��P"`* ���`p����k��rD�Td���s��ޢ�`낗��ۆ8��O�~#2���MQ.z_j�tw͑���?�&�ߺ�A%�J(�u;7�e77������>EL ~�����9M��\�L!Q�������h�e�l��(���B� ��Ge�6.�jtkR'���l\��H"B�۫�P]7yI4��Aa��o�cHxS�D���^7!�Ł��Lm����&r��Y�<�~�BA.�g���畸�W!�tw�p����0�H-�#����|��;�	��y+J�������N�l��e]-�W4�ټ/oLs]9j�V|���}Fpy"k�h�~X�!�W�x�6�C��e�՞S~�@6iO��l�Um�19y~[ݩ�~�>�w�ĝ���G�ͼ�hx�I�v;QBk��$�>�\�cO}r��8�N je�>!��>�,�d-���Z�/v8�����7lQ4�])�Ph˝����rG10/Nq�=��;�'=��%���E��c�Q���%��\3�TW3y�k�	��v~}���.b�7�%6��L�z�Fϧ��FP)�|�9e��A�lE8�����Ӱ�U�^?����e��=�EG��!h1�8 �;]-Oq���\��4�R�I�5�S�s��).@8�c��Ovw��n�����W�;
iT�6.�X���>!��U�*G@ؘ2��ˤ�i㜒���o)sb�lt��nF��a�a���~G�)) ��U��/ A�����˫��~0� �������y��x&H�3v!����$�D�5�W;����v<o�����KKI��S?p��oʢ�F_ I�&}:NNF�d�*ՙ�9p������٧�!
�~���'={�G�����RVJc��1����=�C��ѷ�gb�� �ʽ�V>��5�,�L�9S@u��a�t��P�J�����*�b���?�a�=e��8K��\C�s��]I�I�p�6#;7�����	���:�� ��T�,���o8fI��Ť6S]���HV2���k���ԟ�N52~l�P�*�/ՠ8�w���96;\�~J��N�!A@x���d�@� �ѽw��#�U�`r]��ɛH����|��!�6bo#�|NE�Ql��C���f�_K���i`#(����S��&�b��{�`I� �{hrf�#�r�c�5��KS�q�����9����˩x���U�Y"���T G¾��m��B���s����u��] �9�I�8�N�
Re~@���z%��\ω�H2�g�9�[ ��O5l�������)j(#$`o��i�f�L���yfZ�~�|1XgXV�?�`
_��BZ�D]�0���/54�����N�6ڔ+�I�<��2ﻴt)7�A�̓N��F��9!wO|]j-6��V|/�!�BW�d<y#W� ݓe�י�k0��'j��#+-/�%�Eu悓s�Ʋ�Ryd%�V<8���v� ��=�ȜI�PN9�Og�*kf}���k���q�\&[	�`��VA;�%�;��V�!@}���K��f��u�2 �?�A�2�8����l��}zq����^�;	ś{�k�9Q6hO�B������L��r�=��џ��U7�����I!���M*�s&���=�%c�\��W�!�͛��J��[rb�Xo;B�ciV������7�F3g,�.��ZJ�����m�g|�B�i�C�pB����� @Z�5�{R�#��\���1��nK��]�%ޜ����h�|��-7خ�Vx���"|�j��7�!"�/�e����ڔ��Co�"pT!�_���kN�B��3ϸ}}0�"�m��q.��9�5?^�h�
����;�@�*㧔������k3>>m�K�3W�����$^�̍�����]�$��Kn
6Cޢ+��e�WYr����r�+e���"OQ-��a&�!^>/@����g��:��G�m��h<��y�e��ٌ(��G�ֱ+9�˛ix��9��͘Jo���	��f�MV.�sW�k���:r;�H�zyoz|���L��u��$s�0������?&�f�?��[���F`4���{��T5�4A�6'A,Aa+�v��N.!�w�~��Ȁv՟�h<�N�A��<��}a[T� F�V ���#���:��/�?a]�w�Rv6�>8$9��O9�{A��<K{b���������p��F��r� c��.�c���@
C�Ҍ#��}�׃B���5��)%&�8+�O�����AC?w�Y:fܳ�ࢬ�>�y)Q��Χ*��2i"E��I	f��if���G<�;]��-��T�1����V���u��d��!HqݲE����0a�Z��KU���T����IQ4���k�ĝ-T��N(	ʹ��c���C]a� ����'�DJ���@�8�9�bW��;
��a�&e�E!{���8�R�Ƨؗo]��u��_@݂?��U��1���J�i��3�¤�;�,����v�����6���̐�V�6"�P6�V��y��_�	�#��1��c��h��I;ʰ�+��	���1W���� �h�x��O��=��鑫��0�u������TM�����w�3@�f[凧osX�V��
��X��̤֗���o]Ƒ����UW<��M����I���-�|�k�*��:�ԯy�z�� �G�Wjѝ���e�©B���4-��Y��LyIhH���h�7h�	����g=Ōo���(��ӮY���#��`E����էy՚�����L��Ϟw��j���jS�
8���Mr��+(j�,�{7uW��Y��UX�˕d8��ޭ���>Sr���X����L�g��M#���$[����Aw�||��׊��
�Bi�p	k��B�@���j͠f�&��` �HA�6���M�`���e���&qumɝ!�Wƾy�L��|�������Z�������޹^I��~)"��Y~�fL��H�˙'����1$=�ԍ>��(a�W������E4�I0E�)Ӣ�e���dy��,LŸS�~K����I�e�'>Ke��2�) ��[���6{�5�����
��ϟ��������!�����q]]01Hڑ�\*�gz'�v�`��4�!�pN�_�~�;�5k+�`���W��O8Rs�W|� C�P�p��J�*nC�&}s�h��]P���ٵ�~�{��ѯ�v�?���2�dଶeS8��}��e/f����	���x�Ŕ(��NwΊ�qW����B$f�&�$�7�J*��!9��O����Hd!��iVN�
�œ�)�d���~}�^<X(�w4��2����H��*��I2t�&E��;Yσ6R)���y�~AT��ρI��������@�+���帊yT�����2`t��K��;<���n���U�r��2�[9lxb��D{��������=(�R��a9P�'_lb�܉C�V�e�X
p�:(�_�@���Q���^��ߨw���0܋�'�W G?���;��ZK�n���<0:tV�~�xq�i�
�1ȃ:���e��f����%�������c(F�f��2���b�����H;;�:��M.�X"���݋�̯49��!/��#ڸR�5�E9Z Tt&޳��uZ&[�8E@Yۙ1�7i��Bd�G�vKyNJY?m�2�}�M��d��\�1G_�/�_�3*װx�Eh�����X��(9�������'8��|-b*ɟ#~C:k�~n�	��c���=����S�7im�������C߉�$C�>�� �Mfup!���Q��3�O@t^��릳`�h�WB
*W�τ���㌖��!#�l����-�z��J%��DO]\Y/�h8�7�Ûat���Ɍ ��%���R1��K��o��[�$b+wio�����c�����rjD���2נ�:�%�'�>�>y�����u���8I���: �� >����z0�i/Rt ���ߟ�'n�F�6=N�EK����˄�۰uQ��И���K<�s^��[���H�T$��r=3� ���2�/����ҹ��M�2�Xw<���^`p8�,ˏ��3�!<�%��[��u�FD���XU�
H��Y"�G��4�`﯉b����B�-ݺ�%�嫆m�E�ֲ&� D�adH��f�U�
vԴ��:(?R����P�"a<	S3�J!Jt�kR�n	?��F�B�\T%Nm΋G�%�}<�0Zc3{6��Ϊ�w�Z��R;���dmiH�cj�2���!+Q��'cw�2��߶8�������W;�����IY3�T���E�����&�WNma�Z����2�mҤ�~O���#`�&��Z�����i@�*�iY��69v8u}-SI���q9�W5���g���B5C" p�v�w�#�y�R��)��.�"�X��9AS9+E�'��+���|��HU �Yqi��2�
vI���� �9�#��`�q�ޯ6g|r�My?D�3��c���<� �?�j�A7|2������%~��:����H|)�!�τ�x�'����Yx�ꑆ48�W,W��8�+
�x/�%�`эk]c�c�H�-�,�H0.5�s���5��A�8\N����� �f)�!�Տ���eG�-��u湉���*�ހ�(�r��f:����%[��S���<ī�=�ڡ����nԶ�7=�UsTI���pI�/c$	�o',n����J�p[ތ�����ZL��;�i�V�!W~E��kb`t�	���	LکqS�����������ܚ��	`^�+��e*_�ۈ�2���K]��%c?�W )�U�*Lr����[}�b�{�R��J��L};D�gL�w��}�>��mݛ�P�=2w���LV�L=��;9^�z�l�C)��?��"ٯmu���߻J��Hkæ=-�Rz�6n�`;vl�矧��.���v�fe�]�y3ݧg&6>�+6T����Ee�G��
���@rC�N��K	\���v?�8�ƿ�[O�(�nJM�QP�ͫ��8�z��(�=��%{�\�X#�"�P�l�O���jKR����R��V#����/+W��G�;3#-N+<���"�Y�F���ܭm�yP�i'��P�6���͎�N����H�|n[��Q�N��VH�MB�E�MP(�̭������,����VB�ІYr�.n��M��HߠdbA�pq�*�}���<�������e�s�I��,��j���?����%���W��Vj ��~y�)�v�׭q2��:�M�:C�;�����G�z!��P�H��2�s����v��+�*��C�^-�I_�ŷ���H�N����[���䨘�ݥx�.���� ;s�U1Ι�LW��S���������m�'J�2u�zF[-��Ζ;M��0��de{��%��I�1���7��Hff�����Rj�q��҄��$��,�J�٤� ������	BSCi?�\�6���j�߷k~��S���ʠ���t}KO(�q�xX��-a@���W
ξX�iNq`I$O���h�i@'��v��dðq�Z2Fmc��m�F���6�]� e �"��""�n	�FGJ4�q"`�"*���'��}?�q.�H5_� ���+l|..;��2�1Pa�hdW��R	��Vλw��W�(�_P���f��{H���������H�㝯�������:q�5L��b�۷��C��B }ҭ�~�]�X�-ϕ�F=�yxRENy����d�zgw����Ik$!���BW��aYNI�
����+�L��-ɾ�Oբ����#�����ܓE�4�(���͂��Ɉ�K����.�����'W{����d�ux�{�_�#~۪r����sjʋ/���Q?@�/�N��tB��S���ݼ���Ǵr�� �������+�
����[�o `}���\|2?Ѧ+�n\Ry�������� ���i}Iox=�������V�T}j��+K��ϥ�B;�obw_S�軲Vڦ!+8H��X�K5Q�V��`���C'�)��95,~`\����x[�cND�v����Ae��W_Ç�^Wo���p�@�I�����I�����`vQ/Y�@<m`�����&���I�w'�$��GL������&�����`�:�R�돩��=Du�[l���/b�����'x=��Uَ��v�9����6:��F�T���w�wb�"Ȁ1�OԘ�3�Ėj�o�~*w�t��ՠ]?N��/��Ŕ�_-�#[EݯZ�O�ں��ks�p�1m���Ki��1�#�XKI96��Fw_:��;˅����o�<��%ZP|S���e�J�Y��Pn1��#�f��j����IQ�O`����~�')���/���Y�\��m�=!N!��P��b�dR��r3Q� ������F.�3��FՆo�4{DԴ�"@�X�A��|��Q�AC�#X��ղ�̖:�Na�h���я�"Q�5�}�SW�34Ԝ��8[q9bm4��GDh�m�C{�hE�5VO��*��Y��]ʂQ�6�!�Z�Bj���}��f��p�LP]1r�o�m�ARC���)�ϖL������'�W����2�����E�\�3{�x��q�	
̖xCI�!`ѳl�p���j�@�[n�������5�W-�ߠ ]�j!�����q)��E߷B�8=́O�f�3m��N��Ґ��y��>���{+�-�ߘ����`��U��$\v��B��P�9 �ur<>/PnKd�z`�.0�j��B<�)<O�	KW����&Y:QNW�?a0j]�;a�I�|FLp[:��A���e7����լQk/�Ev-�������O޿��$�ARV[�����>�Oީ��L����}{l���X������bC5���[�����$���N�5�T�` �QX�\�yf�(鍷]:�M.%5\��B���#̅+�28:��8vR2 Ȉ�:Gǹvb ��$�j��.�q��~u��3q���<"�j�\)P�[�pJ��u�u����g��,L�`޴�t��~zkV�/��m�"��KΩ�`�[�[:��z�T�����\��^�����c�%�'/�"���k����|�0м�(�Q�ɷ0���Ŝ��Ǭ��x�D�Iۉ��2���"�KB�X�4"���?�a�d(�s����C���C���������������H-ȗ�
�Fࣁ�����+T!�Ϩ'��%�1U���Z/�ځ�f>��S*���Zȏ��1��߼�M8m�9��o��A$d�2z�AO^�r�tn�ף��i�aFρ<]����sy��E�s[����J,X��@��%8r�K��6�u6�7O"$��bK��~:ؿ�}�ܖd'�:~`㒈g�) ���>�|S8	�<~���YǯaNE�֎<#�h�7�G��I�Ɵ��J�k|Y�ly�: �&#�����?ޢk��}��;�Z��.BH����
E�RS��Z�Ԧt��>V��"��$�(�7�#�#�;/����܂�l�m��-㖓�`�,"�)�J�z��t7/�qzWK�D�+T�ɉ�O��I˧K�O1�)�pM|�o��M2#l^��>o~�!ws�����������;�x�t��GB�8B�>E0�.ְ��U���O�����`�,'礿�V]�}������t��E��#�I�A{4n��eQ�A|!^DlZ"��Ť�u���������H���g��2���i�k���)��S`
�q�?D���a�犀tT�V���ơ'ڄ�4��UJ��5�[����AmPS)�v�P	^m��0�ณ�v�	+��)&�����Z����R��3pL�L�[�AQJ�qr���������e����z4:�P"L�H6؇GX�qa�A?p�[���m�8�m,�z�Go��+�<fGX�|�[[%o޷7��� �FELַ�U��ȯ�D�I&x :����|���E".����|q���)���>[��D�DVf�+J,����-.wA�P��w7O��i:���*3&�9B��Y�ze4��z�X}�Sz=��/]ڠ̍���꧳�}<�����TO%��7;��g��c�� ����gRn�7^�2������w�L��,��<�����%-	�>
O�0H(�r������������ۍ~p��na��4{e�|��"B�g;���R���"���.�^c��D>�P�������(��w�NV�m^�?�ʼM>�t�v�u@?��#w9[N�g�W�85}Q���a(a�cL.�M�U,��[ر�C��w@ޢ��q�,��1-+(��1_��/ϯ��07��s�kMmA�
�xfTm�{8z����E��>���wD:�H��͘����ȑ��7�hH�r� �|��	�,��#������t'<"4�jk����+z�`~����Y]d�2B��A������~J�+-�Z-"��R�U��^V"���C�SqZ��v��7PI)z5���C�Tַ�����=b�����0��{j��H:̭זs���P)�}n�����|��HۣaNR�r��vW}{� �%��gm���G��
�Fl��HK��?L ��h��u�3X�2�V=�T[��Z�4eY>�"�x�Q���U �����^8���������7v��'��u8�B�������#uR�m�&+U���Ҡ�xJ�3s��8��?$'U�9���`�7%�&���d�w_�T(`��yf��w���ބ��B��V̳(�7�ý�.y�獚��a���]4���O�k#��d�q�ի>¾+�I����˯p4�����Ţ4r���秲�_���L�ٺ�}�_,�ޱ�d���N�#�	�z�M�� ����f|'�Y��ވ�!Wb�8>���a"�Y�l�{ꡔ�!Nq���7�aP�pgWS��r���hǾ]��2)P*t/b�N)����3<z�=J	B�jB�T"����d����\���4��	���2	I���.녉��05���G�eA[{���ǆZ�3Ģ�!v��B����a�X(�(D@we)(v��>�vp!�HY"�C�L}�D��b\M���������S��`m�k�EUg��A�Pw|��A.���6-`-c�s��X����CX�J�D�9�5�����̷�E�*T ���� ���[�F��'2��4	s��!)/rU՞�U�f��]��=���
���X'1��{�=rN���b�Yʀ��K^�<\���ih�g&'$;@�ĳ�lq�F�D�қX�a-�j c�l��+��"K�/��E�R���*�!^����f��n$��</qa�����r�Zh��)]��X��:�jx����ó����h|�5 �7���Nফ�}�A�F��x�OW2(�V�W�ޣ�?���O���OK8?r�_�5I�3@:��[)G$7��T6p$��ӭ�c[BY��c�@w��@MQ��	;߅Y*Ym�ȩ}���F��su�g�����D'Y���I��C d�׵����y�+V� Y��j`���_'29�Ǳ�\7��m��yf���
��"x�MR�:���Z����[2��x�g�U�m�eZ�B����������@�ս��}Ġ[����˝�p��������,(�-v���o�0R������S��4��x��P&�?U�(�]=XʪGf�Dr��D����V��*4B;H���~�E�ӻO��25������?ȍ���'�);���CA5�	�f �����VE��t5����C��P� 9v�R���?@uW��x��8�%�?@2w��l,w��0��c�2���j0��������s��8<)l������^Xo'�^�5EDH�3��^ ������늑Z^F�^��Q������<mL��������}uf���v�o��av4 �NMz���Y"
Vj�%�z����Z�������'�������P)K��2�U��n��o���M���j!#�N;��F9�+[�ޛU��w@�ey}La*�Nˢ�w�H*�)�LB����Ε�)f��h4��N�^�R^F�6��Ӝ�q ����C��ǂ�F�1WϾ<��u<��-&�&�Y�嘠P�Ϭ�\�][�]���:�3��i�{ �@Y!�*�(|�
�{Xy��mC��1�M4�*G[WC�mMH�;~���7oI�^�j�Vy?��&�W4�m{%�h���E�#r�̭�(�j� (����;V��Ù�/�6!�^{z�=�e�9�݃�Ų����6�5u��Z��#`}��ϙ��a���PdG�[1a�mw����+�Ц��m��B��1�m�f�fI����Le�h��8�	V�F�]W�e�<�yWcIx�:"܌�(|M)��8.t�Q��0R%�Ɖ
��y���xt҆��\��)��e�7탮�A��Ȥ��ŋ�Ji�0۟��������\�sҗ���,2�����#��ש(�{+f��WG�����Pq�kT�#iɬ�$�&4�8~���T�m9%�^��PR��<t#ZN-�?���D=kPT=�c��V4�7anjeʩ�E}�t��N�IQ�us*t~��8���0�v<i��������3r_H�
#���%e@�u�l�W���q'���q΍�f93��*Ҫ"��Y*��S��xɀu�*�|��R~
����+�3s��-�_bbDVR�&��W���@��M�c [��*�%�A8��T���5�ƗU��`s2�K>��KV�ᰢG����(U3����#�f��v����p�&$<M�v��ѭ6+�~�ĐGS�`mz'�_^A/Ga8n�~۳ؔ�{��j�R�O P!<u�`�_楐?0;��h�����D������D��^�;u����jE�T�UE%��m�/�`X�5NKJNg�p�?����b����^�/u�^6l�?�������B��L:�L����X��Y~	�~��?r������y��r�������7<st��~�k���rD@�s��:,$��=h�5��ѐ�JP��Ȳ}�����W<v�Up;,x�~�?�;4�S��J�ą�}�_�׀�����$�f��\����O�jB���d�;M�����1�!�S�orR��O�6~�zB�"U��{y0G.4Ě�.��t�%�JpE��XHO�@e�$ޏS�S�S�q�p����l�~D�BF�x��)�mGC�rMb%��R�XI������8�Y�U<�Z��u 43;��2X�e�&WO��ȝ���9�U
�u�
�����s�� 1��u�uTC0G�����H�Uy��N�[�M1���=�T��fcټ��Gr��S�Ls��bfo�i+��1^��c�'+�MR�|��Q��}�W�G����=�'��{�Br���� � _;��	��su���h�|C!D���u*��5X/�y�Ų|�G�Ǻ�a�m�>Nn5����[�iC�QK�.�aΆ��:��[�i,��Gj`�PI�nAVM�W��� �%yRj$����}0����qr���'P���Л'�����+1�,����t�H�V:��Dur��{�Z���}0n�o2�P�*0<��$c.8����<f�&Q)�Lg�C�@�J�	@�E�r"����tKX֑��ᮜ�8�,A�|-�&D��xaP��I��Uţ;�7H�I/(/`�\$��\[�ߗx^#Y-/E c���z�Z3� �2S3�;�wF�)��i#T˝�k\��Ć�N�gh�)AS��5T�d�ڐ��% V�_/>Iz��w���`���أ�UH���ε��ˁ`>3��� ���0k�*9T������Jv�*#�/r@�����O����0AN� �����4`�D����u���ܟJ��>;<�\���#p7!]�V�6�u�a�"�]sD�5�`D��m�UcDn��I���j?�;R����z���#%��N��20��a��d�1@���3ruM�D�����Ǒ�-�)��Ҡ'�������ɧ*\>ȶ�����r%G��?T[�w�e�]}�N�����^4.���&��	<ޓ_�	*�P�\��1DpX������d��� ��f���_>ۋL��ľ>I)g�\� ����Q|��y��w��e�i�87��]����rL;��:��j��v��K�z��˦�y��Հ���B0Ki�`6�(��?3ԣ���,��4�
�gT�̮^ےSd�d�$z�9@�A@6�zWQL���Şޑt�K�H��(J�cF��t�A8eV�5�`H�\����eI�n�Р
U7��g�Oo%9�/�*�0�f�����	�d�|v`��G�A�[S��)R��LlPF�:��d�~�H`�q�%̈ytXڹ���F�����j3ٿ�xpK�.$����y�E�s����V����,[����*qb ��kJ6��t�#���[��6}���o�~�D	ѵX� �#ֱ/�% oHC�&|�>&����5�"o���" �	�|�T�:�h,V��h�s���77��{� �o/5f��JMO׼��#� �#��Rn���UNK�`/�9�M�#"f�t��>�.��ބil�-$5{�{�0w/<�����$�`/�q�C�L�:��\W(7!T��￼��5��r��\�xn�
\��k���t_|�vg�� ����޴5s���̥�J[��<���%Ҡ��_�M�D�7��6N��lQR�]UN%k�`γL�:���"a�nN�V�����^���_��?ls[�~����_�ࢗt��`]Vݐ+�����;S��B��Ք��6�cīՋ1�N�l�m��!W�>��%snz������ץ���ď��Iuz����(�c ����d��@g�6�<F��oz+�zN5$�]q9����y��į�f��Y�������Bʡ+����>��.(��oV̯��<z��]���v��ó�OYʄ4���)L�2Y��uL��>��qJ�v��
JZ36J`�R8/�kv���� G	��0��H��/���>/e����-��+$��7V�W�B�^�\̏z���MqX���qlH�������B�d+�< �K ��[�Z���� ]�i3�֧�d�܉&Q�dP�:�)���B�K<���Rv��G1���i��䏤�H
� 7�,�_�4X�\�������5Q�LK|�X����V�轎�QI���5��l&�{����̫�e��j���E_2w7��p��)��f�y=|��.b|���eL�HB�������R~��-.R�7�n��)$x�Y��IM�Z�j�e�8�fx~��4?W����J�����N:���DܣU��!��:�֞��g�G��!X�	�YuO2����F&�� �un�ge����NW���y5{B�h����:�ΠU�'(#39�����D:`	�n[��u8WT�5�2^I��^�	N�l�p��e}P���,��D�X����Dd�-$
���E8�W%�q��B���s���L�?.{{���i�wO��P'����d����Md�>��i�.�ѡb��c��1�Zxoa����x�6m.<S7X��q�y��q�[���3�\���	1!S��a�t�\�m��299�-��2�����7���^�+�*J7CH�3��{��o4��2j������	�����z�>P �r(󾸅�7a�� Ѽ��{�=�b�s������Ϥ!*�2�ʬ1M^)���0����B�T�z�� u��	g��a���ñ6!"��Z���]\|� 3���̢�d~���&*��W��0��ǭ
�F*aso1.W20J�^`���N�%����4��·���j��h�����Yʻ3a$W�_ju�z�y���	�Z0M��_��UKW�Uk���3�cy��-�y%�ɑ�2��gd�5*w:X�E�NRṇw��3��b�ۊ8"�?S5c^���͛FGز��d�]db��)���c��Wޔ�o�W�er�"ߞjYwk�'�\R�͠7=�W� �����T����[�7�������Y��u�j��?z�U$h�&c+am� ����^���=_����%ڼ��,#�I���Yj,�	oE�<S�t�v�J�^Q���5b��\y��iBoPKg�h}$=�ʙ�������bc����sQ ��z#�I�2�Z`X��x���Bf0��g�֧�(��f���G�n���#��yr:�P�N�#_�T��o;�����.{�a\�ֈF:$AE�S�2�6J���
�~����uN��UDb���[e�B	����7g�[�aN��~�_v�<�쵿=����;�Э��͐���1g�����W=c�����}�js��X�OZ�q���w��E�W;��+?zI�L�4��jѼ/�󠉎�iũr�O��iԠ�
��9�k %�-�&�����0�(hЄ��>w��f�4�w�v���C��~zE��3��M�����ǧ9I�2roM{e�>��'+y�a��⚹���J�ō�2K����c��7��M����+���nh�!���h�P)���P�����<�2V��}���X�0��N������+1>L��j�<�����o�a��p�x/�W5��ud� ��tSz�����]�����^�g� ��@w	��N�e�c��zuc^F-5�Y���6����R䉛�*���WĈ u��/�T�t��;�&���<�v�ڻ	R/J��|Kb=�P�L��B�f�Y���&bQ�I�u�N��R*.T	�b X�3+������	�o�Z��"#L���?5�K��z�h|)N8T�ن��Ď�=�o��Z�X>'�/����#�I�	.\;��G�?���L�7�����y?~�T���scQt��7�k���\<���.�H!����E�n3��bˠJgTU��<<��k���Rv�*_r��m��."$��/���WS?����ѳuQ�F]:��b�-��t n:���?z���UM����}�G���=	����i[>�4 "�G ����OF_�g��w����ћ�/��?2@��r�	=G;Q �T�<�N�С��Es'+�4vJ�kg[�ޏ�89��[a��h	s7Q��K}��վϕ�=�n]�t��3>Mr�71����-x�(��U���MC��{�i}}f6�烫�s�֘�P�pr�尩��L�������)�g��N <{<�fy�����(q�����/�G`0������?w-�^�<S�6�ם�:�	9����E�����x}�J'�2I���1t�{��1S����;�������_W�8�h��msA��2��K�Wu*��A:}a�%�W�o�p��Y�4C�%~!9>Ux���v�|�J����$f���j�x;��{�@˪���,�1�rg�Q�����a��ľ�|�a_���p�"ᇼ��O����9���S�W�Iٹ�wp��3��䂔��@��D��p�U�)����Br���B���7�wtx_�$@Ɋ�ю�z��8�9���;֟�ԦZ��U]B�y�v�Qr��_v����t��H�d�O��:RW/�v��)"zJ	��D���Qh�bY�uX.��"���lnuոx�2w��yR&�o���C<"�}�O���&T�}W�FA4S�}��2ZU{���Щ�`
q�"���@sP �#\g�u����#z�fX�hr;*��0D�򲹸G�5���G����(,2�P0�B8�&�+0)��������Z��D;c��2����*�n4~l�Re�U<��Y<�Qe>Ͱ�*.?��Be ����q���f~=׊�R��&��!^R�5�.L�'�| �v��p���n�ځ�@i�V�KQ��AY}��@��2\K����j��o �i��9��4ƾ#�>دh)����&����Kn�%�qu;'q$Y�:�1��پ}�
z�W�@��ŭ�Q�Q_ޗJ��\�@�/i�6���KZ���"�3E���J �v4����j�ρN9�]�+��&&�����S���嗪^9i<�T��ח?�>L�0��t�A/8vP4Fx�Tp����G������_�?�աW�D���G���O#,��*�k��kHb����n������e��m������v7��h����yԟ��RV��9;��E��s�qtL=`�(�
ƶ�b�k��r������n?��Eݚ}�ͳ$4v.��s,��N�4
�<N�s����,��D�(-����f?}�k:�&rA����_/�zn�8��\v�:	��`�r6s�0��<W��'l����u��{�^=�a7�"Z�q'%�?W���A��-b�I����/����)v�8@xi�/���Y�(��,�n�>�=�"���?���
鳭��>��U��B��ra�a3�ζB�����/��>��$�|/����Pl�B{ޯ]8j9Y�ۑ��a>�|\��Q�{@�\}��g��m��?��`� j�7x��j�������u��kj��"��V���3�+�a7_�3��;X�j�gq�n�DɐI(^�*�aJ�~�(H�x��������Nd?��(�n���$�*�O7��:ə����<9��p�3n��pT]�˴����rܻSt��Ɛr�A�z�[��I��g34k[_�tfxC��	{'�J�F�S��F�#('ٴ?(����u�����˳�� ��->z�3�Ǚbþ�[��@qUp�������R ��m���]������d�ƾ����i�py�m�&�������N�ۋ-Y��ea�6h���v羪 D=`l�﨣t̕}s��$EG�My� >�vW�DOO��H��~.V�!^�+�Zbw�����c��Ί�XB(֯L��%��XF�S.���uF��j%$����L;�C~��yA���H�F:�i�i�<j+��&�ħx���f�4~(e��)�IWU%�Col���F�Ť�0�.SDԾ98C�Xg��1W�!]yXZ(t%*X�ixa�Jf3P�bI#�&��S_C�;]so�?�`=$,���ce~���հ���ґ�m�'�+�c�a�O��w�Gǩ����A#Π�2�=Ko�0z�7�Gi^{��F|�µ�g�[l�F��=��?�Ý&�8�푧|�3�(9��a�M�6a�0��ѷS��7�P��4z�]a<pzj�.=���E$���`(�|綍���=k��ț�}|&��Vո���ZQXݫ	�T�຅��v��^.8����->�M�n�?�b�5�_H9g��Z'J�o��õ���+�����srK�Q��3�C o���_�"�z�q�lV:�ӷo��̬���<�uk8`�:[e!��~C�}�6͗,��[�Zb\4-�R�����K�E\�ސ4"UR�i��֔�f�tAL���[� L�(�;������x�9�Ǯ
���yC�8Kw��e����9,����i����c�^��C�Zj��\h/邎�s/ؤ[N����"߀�N%�z[�q���[?\j��T
�Z&�D��$�JY�A�B��bC�ļU���:xn�,�)�|�m!�8�
��;��
��|FU� Sn���� ����׎q�D�/�HUܞ��v݇��t��Sp��)QO�\����_lu��?-N�5�����UGfVP�^g�Ϲg��ƨC�H��AB�+mT�^3���s�1��ꩂxG #~9ʇ(����~�=n-��_��>�F��2�?�6␂�$���g-]6[r̛E�j����nhe����H�-��G�rl���S��~�(2uX��j�<N����&e�k����pN/,�b�AJ�0o�E"�y��[a�V�����
5~��=��j<�Y�8"�C�&�p�[��ʭc�)�h' 5�K�<�r�%��{�5�X�3��}�Ry�����6��n�-?��;���'N��r��NS�1l��?E��.��3ǭv��mS�ĥ��+���$��,�5���SLmFf+�R"�2��h��gkӑ��>V�},N��*�f=���l�UxcN��A����5������q���mr�"����Π�)СY�I��/�i�;	��?ڗσm"Y3�����)����:�����Ȑ��&C�2�J�UH0���q&��2y�,��z``�xن�M��E6W��k+҅&[��7P��[	��d��}������Չ��ɤ�#�|���`�`��X.2IV�����)q���p�誉ذZ\:�W؀���z*a@)S�3~��ө�VR-���_&^B�����[:|&M�|��0�ږ����nx�cm,�K)Ω���ٺ�/�a�
m�!#_4!&)]F�uXfԾ�M��O�[q*d1"d,JqT�}T	�wݍXIE� H�Cp��Ԓ�Pr���S��b��$ЫPkP�c��Cʙ$�����R��S?Zt�LF���]u���ݨw�k�du2��8^�*���^`3�l�2����N�?^<��?9���h�'3����:j��>��6��!c[r�V�St���m��iױ�L\�Ϛf�?�<0�A]p����B�W^`K������n�8H�)w_�@��)eGt^�2^�o�;�� ���!�ʦ�#��/sm��`�x����p2����V��ʋ��[��W5O�`b.ym��(?Շ �-U��z�*�?�?�Kl���x稢	N�4�]��;�f)Fի6�X��#})�^���H�c	̰���=[��B����;;3Y�.���
nL7u6�;F�&��7;HE��=�G+X������p������4�E���26zXjv������-5#�3������ر�w�/��=��
JU�@w�;m�[op�C��Ñ5��:���j�~x�j�+�lNx�6m�_\��1�`ʈ5F� ��c��������n�A�{�H�6�	-�����u����:O�K�U�ª�J��n|Z�@���w�Y:£����H4�uBF#l��9�%���88������_��ԼV=\�#�I��2��!�-� �V�z�gy��燎��\Ǧi"� �T|������P�ۗ+U��}�twT�����喳�E�0�n	��Y^o��[a?��8�H��}6n7Q��Bx%�]�_3/̱���v�B+�}�D��ڂ�/�cV��_���$ݸG�Ĵ�y�P���Aĝ�N��i��j	k��k#B�4
�����;㔎����r��޹�2��wk���5A�ʹs8Oy��`�E|�\�Kv��w���g���C�2�YAny�T��9� �9��AIvIѲ��9F��̷�Y?5�	�Ө�~-C�iQqb�"n��l��;8):����&�Z6+Q94Qϧ�����C��ۮ��j\tg�CQ���>�F�`3�
�H�\JڙE���E����,`(`�6�ُ, �NQ�G�6(�Z\IྔsÚ�X^�
���r�i-O��ş�Rﱇ
c�{�[�ߣX?�1Ŀ���~*l췦K��|'>)��4��8��'ե̢���c�uYy��(������F�x�6�cO7^ě�Y��Q�OO[�ɷ��wd�	��1"�<���?��KV���J�iY�����N�+S���jͲ��O�49f�!,s���s��˔{s.�׵�F	�������
z���AwJ��?��Q��~G�Z�.�G���kⱅ�%��
���:� ��L�o�!�������u�i<d��u��-����A��H�3-9��JE���s�K��-���Oy��.�~6��c���&��6	����W�&�[��*ha�j����Cf�R�=�E������đd�JI�i!#[��[�g��C��w��sL�^|Y��Bl�J�Ih�/X4ocZiV�޵
��?�/��4k{���
m\��wZK��or����vo�����+iڹ�˿�\�x�Ჾ�xo�[�!�aP	׽�*@DB����aO����B'�ꞔ���}�\���H@�6�E�����7��O*��ԆS�?��Y�VB0��i��r��k]g�K/ �c/Q>����6���J٣� ��Л���QX;���=��~!��)��a���I�7͵I�⽇2+��е�� �l���Z0����z²A!�᯴�"��G�yg�&-�j���g�>s��9ޚ�doV �m��e��GmQ��׵�=���A��JG���Yń���]$�
�����5�Qpn(
k�]SZ�[ڄSr�醴O�]ts<���}K�N�JJr�cdN"N�nW�N>��]$T�������~W2Ԥ#7�:3�沒]���g,D@�9�����tF��`����n����b�
ѻC���̯q���V���␤���҆"�u ��cي���3�gq0�S�X!0��Ϯ\��;6�@�*�I��MOi��4IU����g2��?���DaK�M�W�A�Ӱr�E�m��}H���O�{d�o��^�6���u*6��>5g,�%C�'.Oؗs����d�:G�Q��#�q$�`����0��bS?���0c�,
�*!���'��+��5�����"�|"���r9��;����[ O ����7�Lw՟�߫*��?\���2���>�V�Լ9E,;�I���I'�lJK�x��o�(?�|�=dj�݁�XA�;,�<WU���� EV�����[ۓ*��E�s�@�S\�2���u[���/�n3��������W^����鑛�E:��k���a����{[7\<���op<������;6�kӶ��y��ǫ�}.5��Q��j�g��=KFq�n"�R �5Y�b�Z�AH�Y_o�0��)i72��Ut��T<�G��Wkn�rh�S��ֳ�8/��4�p�A}��'��eH�f<�|Բ�����Z�9�Z6db[�@{��ꭹ�o���h�~�cH&�Uȟ���KI��uкBj���H;�ս]	�e�������n�r�C����p�Qp���钙�@/�hx�Z�0��~[&�%XϯqD�#c��#I������Զ#z�)�@Ie�XS�S��d����;��!3�A��7��>�T�����Q >������@�"�vBq)�w�S]���$苄 [9f��ƈ¬���Ȗ�l=\�W��[})+��5Ц@���-�aۨA�e�0�yͤ\e�?����WfIά?P*�x:5��D.����8�e4-d��{�gFtAC`,��<Sق4�o*����u�����X��^����l	�z�ኮ�sw��c*F,����ފ?�����_� ���>RP�D&8���K�?�"��/�MR��^�z`�W��
y_�����=ele��<�U� ���F�g�nA�(U��y)�'�������#�?lT)�E䆲@`�Q����$Vd�ci�K@�S����֦���?�厡�p�)�)�^���>����U%�R�r7i�S����Y���SZs�]�&�>�CC_Q��ی׈¥DTD��)�ê��w�N��G(U��p�U�N*�性����HN�qr$�>1j}��ڭ�SB
+l��=/a]q��J �+�6N��-b�Y��w�*��F�e���p%|��Anp�����w��P�H�>ƨ
 �k�h�*�F�,�Z�(�d�Mj-T=t%9����U�]����.�x��w1s͌��f��N��șmnQ,
�$�R�3Gs������Jn��$�%~��?�߯���4)9&�R,�"�ej�#s7C�"9��9��oƌ���ߞ&)�mA�\��hK8<�,�@�P�mB`PȀ�g��iɴ4t�`��$d��K����P�C��|:m�
�k�e�᝸�t@
ln�ԓ�dF�cl�k���I7C1=3��C�\Q��,�g���V��!��P˦�&wx�9]��z<���;M��j��u��=�J��~[ֺC�kf)OVf����L1���Pw�e<G�>k����6o��q-z�Sy�����|�����[�SF9��>��M�9�9��@�D&�|Bn r:�Y�+���O�)n���Ze[��BhJ�~��~+����.��Q�D�Yg��A���6+:7/��X�������;�o��d�h��m�Z��Z�$���]��LԶ�35T�k�{R��I�kR�����&���w��������dp��4v�G:�GI4��7����S�x��� YU�U�»���<ߌ&�9���D�VD�d��<�4�;VOݲ�,:�lX8jbb'Z���y֍: �k��tD�]O��>�/���،�Q���;��bZo���v �Y�<��{�4CO����t(0��%�&��?
����`�	�틕�w�0N������ϴd��k3��c�w��4�ʩ�~�x5U�+�4�J�Q�ܒ�'�I=r׆=�»�67��ޙ���@J��}�iukM���8�E1���M��q%�v��� ���|�G����v�AT0򗜽�)�jl`+��� 5gRa�kp���IO�P�ː�/��|�V ��\��p��(9�����Kj(�u"��/z2M+BP��Q)Y�I���!y�블,�a+Z/�Eϥ?��2S�/@����Z�:",�ȱ^O�����d4�S{�p����HU��FF-h\�֖�t�h 0�"B���G�c"(J��2��`_�UB�>l>�qD�|� "�Bm1�M�Xpv[��U����i�N'�$H8��t=��I���`04���M���,#(��e	Đo�N���j����)h@�����0 ����z-��KZ#}�Kځ鱰Y������$l���SL���v,���С
�[`C{=#/X���¦��m1��8=��8��c�nJ-�)��0�&}*-�0�#��%���P�5.��ev%Q�ۤ�����x=Ȉ�P��=#%��$#����-Zv��m�u{�n��G�+�>h7��b��?3R��ᴇ���/6M��6�_N�2�6�3�߱�u�'l������'���{����ܧմfz���K�<�t��+Lj��Y��̈́8�O�B^�f)Eh�|I5;�G0�T��uL!jTnU��N~k��ux���=kZ7�A5��1���UG�ω%���B���J�\���+�6�[�nY>�:�K�?р�W=�b�����Wǫ��8m���:��O|�2�%P>��� �/���:zQ�P�� �ɔu	�p�Ù6#�Gm���f�_��%f��l�tc���6�K�.��ސ�乶}D�S�����r�Y�ա0��3�57�#t����=�r-���g�t/�_6�m�w���ry�Q�R�"����)n��(�6��5(cK��W'9�G��3��8ẕ*�Ygl\��d�l/w��fX;��i��Cށ�v��~�/�����ݍ�,�~��F9r6r�� u��~[�|�/dsݲ vd[o���xA��!��?]����?��G
� [hPt�86��lvb�a�'���?�1<J,\
-��^��g�D��f_AF0#~ј���OO=���+���}��v�Eh�ܧA�ᩝ0��R0{!��ƙC1���
/�9H]�VTx|�4�^-~�����n.�~w>j��J��*&>�}�
��]�rS_]8�õS�?0����NX�Tш�5OA��g�}�H�J�ݐl�������7��?^��	�.z
t������P��{�P�
}!�h@k�%y=�<%����)�Tӈ�z��sΖ������	�������g�S�$��wܿ5�x�
<�
�㭆v_=j1���������D-D���</�/n���{��9��ST�M�:㸷�hvJ��ǿ���^�f&�84׮w}��$[�$9�!����%�0n�Cu�ݎ��A|_��.���M����h�n-����ޅ�w*`�z/�����٩��H��N�:D��~� 70�"�
/�i&߻��<�!k�t��/M�t���=T��1YW��~!V�e,�������<x��1��E��`����bf��6�P��s\2��A~c����vd8��׶Ѫ��wvxn�NI���$�{]��ϖ�m˸����� ��Y~����4ۈ30qZ0�!e��#����3 �		wԖ���RD9�|.@�f"?R��&�HA��d��
l|��
5Z�#]�9�����7��+�N�ᖴ�l�v���H�s���>{0o�Cs�����gt�x���4vx6�
�D|��2d���Mk�� JB�%}j�%Q������4ZsCsŊW��vA��nql\��>���`Ld�y֑��&�_R+������WHM�rZ�i� �)���*��_���l��s%�z��*�WN�[����6�����=�.�l����/�:a���r�'ۊ@�9��C���l���i���K���b��^�lO���V�� XR۵��ib)�2Z���i�]p��N^�k��\bJ�����|K�Y�������\�GR��q&JҋEV�4��FN��b�1c���r���>	�ڏ������3����yg<EL�1څ�غ�X��7����:��5�s2���K]ǌ�x��{^������W�zi^��Q�2��(�Ǘ�R%�"p�ቡS�\)���T�cP���mh'F�"�D��:Vu�����v1��ʷ�,�KƁIȲ���T~�r`hCxL0�\��4��	%A2`j���娀c��A7ݔ/4�5p�ީ��k�d�8D���������Œ�J.�V�����kҴ�����p�`p��h�+B���f�Ty�8���`��׭�	H��c@����[^��R���@(�K]Q+J��T��u�d�����@G!+��������O�&�B��&�k(Yϔn�s� @�>���������	VuU�[�͵4�JP`7����9F s?R�V�:h� t�e�wH�%�s3��6�ׯEρ��h��w��T�H���jk;��s!�]��/�O�I�9h�q�-I���DJ�S~6�ۅL�a��?�Mm��%G`����RN,�\��B�������-!/�'���Ұ�)��Lrtk������T^�!��q#�`f����F��ϲ�f�l������y���!�Z�����'���A��
���{����4�u���Ɣ��H���u�q
�4Jp�����ydQ�}Y<��u�\E�3����rʄ̘�0�uT"K�fq��z�W�����T/qO���X�K��#*2��,�Fǜ�Ե##��v�W8��>�,D�J{�mi̂w]''�����b<׵�$�Le�MﴁY����!,-����n����<����!-�0��S�d���4ᵓPt�zH�(O���.���GG����e��p�4aq����!$p�}6������nZ�Fr��=��-�#�6[h��T��<%�K\j�ڍ	�v0<�xb�k�\��Q�`3B�}�p�~��}�6 �����!ϳ�'���}c���.OB��9
�-�M<���=�d�Yz���,�*�Jյ�J�n�&S �orqf��3}n����Q�KOXU[d��|�xI]��!�Cv��)}���a�S����8 wug�~E�+?/��qD�1x�Ӽzq�8r�v��O�]�;J��8�<U����]K&�)T��K�
1��l�~j Z����m�Gy�O��S���n=񎇒5�_䣝1�!�Y�\���|��~�C�E�@������+�vF]w<�m����}�>lܛq�z.����Eޏ�LSEnHL:�k�X���M	�L���}�!`v�JGO�)k�#fu�٠\�r����1�� �$���l4�#\�����k���:��@��S��\���q�~ϗ0�V�cK�c�������0t�3.\�9�[�>�q��u .��M�����V��9;j�6Ygk�UW�KW���"���J�Ī�<7�|�	���N��Nѐ�F�#�i�[�K:��j	���9����r�2�/��y7�� �����T��M%8��}��'�>zd�*��>u������A�)`֘s�^·,�ǳ���#~u�E$�ɏ��&�T;nT�RB��4&(���M������x����(�J� CGI�B��<�a�T�ah�z�w�i?|��<9�a�����&]�'��F5b�vu�Pս*'})�A8�����p&�������[�j���y+��6��Gܻن�t�^��]�o:�)J�
R���DSeN�^��GW1��?�^CV������-�pR���߿wV���~"`O��U٠&�1�b����Ȼ��u�CJ΃�ϯ�7����zW8���Y��ZU�����\�K�N8 0P��k�C{'Y9|�v�g$���~����^o�� ܈IOO��#���[��5�ԁ�#��M*}Ҽ�T��:-Ո��d����)��wLw�[�z�@OƑ4����S�?� �0ɻ'E�ݷsl)��N����qs�C�ɸ����������m ���#������O��Vz}JK����)���:yR�ǀ���z�yO���Q�+����$��u��|�gꈞш�5!.����p��ueN3(�ޚ�ݡ-�3�8ػV���j�A�]t
Z�R��{Mޖ:&�IWT\��X�1���G%���c�s��|�ʌ��h�����"�C�H��UK�ꇪ�TS_VtN1���q��)d��@`9%��Y�f����>���� 6��7a�:�q�L�Dr�=HO�(�����'�-��R�����<d?s���~M	eA����-�Y*�Nvu�6Hy���|DV c�UoI������w�U�В~FQ�>fq��dT<bG%�*qa0#�B��
�`w�.�cF�1D+^����޵;�5���{ꤒ
�O�A�S#7���� l�E�����{��^�j4Jޏ����V����=Ɉ[޹���~���.�!�s�a=��^�>5/��@fd�G}h��cl���Og�.n�&,�C�� �H�����a2�x�|]S!��!$�ni�1��>�N�8�Lb��%��'!���ѝ,��t!�+a�jt?4��A;�w���WF�@e*��Y�t3�'�@���.�;�B��:���BOJI�R&�A�LY՜ݪm�h���|65l�O��lS��.%BpNξ3���C��ٜ��:���5N 1���m]�G��J�?)/��d�ugΧ� �H�E՝Ha!F��c�x>��}��YS��|i��x}��j'�|��*�5�:Vu1�����FXhƸi�_�;���|�>ٵ��8��B�jh��RDCL�M���֙�´�u>���Ç�J���*E٠ .e���˕R���̴Y���S��{u���|���[3�6+�t?�vM��ۑ�^!��z�]�ᒔ�<�؇H������w����ټgU��}��2�L.�LK���I5��7��}p��^Q�_2�����<)�-`[�ma_|hY�e��;q�ԧܸ8����y��Ԍ`r~�'h�>PҨj2�z�6�C��k&�AWS�g�K�ZM��gV�� �� �5QP�'��6���@�� 1�A�������'iֳ�o� ���
�!&�ɧ6�S�m�$�s.��ap�@b�ct�:/�l$�i퀱�,�+]&�K���uxc�MWR��4��Z@Wp�O�LI�l��TS�&�/���u�dݎ<��آ�0��6�o9��u'օ�#a�� :��qEQ�˗� @�;JKu:W?\��ó?ܦU��I�q��l_%��~�P��|�9���P�P���]�`�����e��Ujʹ�]�=Lԩ�������厂�u���j�(�ݽ�G��d��*�aP�6���)�7�4;�u0���;�Z�l�U`*a}�V��Q����N���{ҏ�a9-מ����V��|��=u�[��ٗ]Z{xR5$��Zc¯PvsIrk�%%9=3v�}6���P�!�d�U�D2�R*i�} �P��&��`��o ��oo<Ux��=�P��kػ�^3�����qY�
�#G��;rĵ�m��nbrv@�T���Y0�rDZ8���4TR��x�iȑ�'�Χ�m�ޟ�6k��Cq����7� 	�?�"�>!U�WvY���YkOeI�A��&iIjI����2ߞQ��A&�iß)iQ:�!~�K���H�	LQg���NM/A�DN��}]lb:����[����G�#���4����\�FI�kh*��f���r�%k"�O�*}`A��u��@�+zS��@H����T����,�M�9ջ�^=�%���5X�[U������ୗ�5�.�6�{1b�����"���+�A�������m^���ί
��lAXR���N�_��cO����_7����m����p�r������H�$ 6��N_��8����sAމ�����/�zd��-:@��}�?�R��Ɍh���Cd�:5+��d������"�N�8�7w���M�%�6�P�J�_͕cSo�;��z�o� ��Ǎ5J%`'�ű����{�6���7����B���	iPs���;��@�<DE���o7�.zA�Т`��<�^uX��zn�S�qƹɂ#�/S^��iY�?J�~B�<��l���,�P}e���͔Ѭ30M�?�	���ˀ��
��A�G���Y�T��me^��ܮ|�a�i'�/�a�<N���2s��G$%Sk����� %����n�{ׇD/�O;vZ֖-��!����`��H�=�L���s������{BUA��e�����Z����rjkx�az��\)rP��=uSa�0Ӑ��Vq����^;�nƼG)��V�����B�/��o�R7��m>�N�r*�s��L�?���[�Ƥss��kbく��.`Z�=�^9�h0��סf���l���8=�e���\\t�j�Ί"�/z]Q�ޏ�LX�	^��hfT����5��`1���T��<�R?8)}�<t��'[Kp�0�N�x���J����6Rɏ��j�K�ݯ�A�����\�Y�?�T�5P׾Ibc(��(M��þ�>Utfw�i�v��i���H�ʴŭ�[�t�Fa�)H�8�C����85/�ʴHڢ�8�0�P(wU5M��}N�9'���ځO�W��y�T�Z�п�sͯ�n�|���f [��P�r��*�����E��u��R�OZ��Is�JK�糜o?w�U���)����B3�vY�%�U����h	��4^Z�Ғ�1_�+b/��\���.��l�z��	�\�ϓ -V��O�8�a�o�g��]l��&ėU������U��B�﨩�������Rs�1v�neD�y��G�GEtY���9T]��| �}��ܙ;_�Ow���x5�=!�J-L�P�w�H�J�q"�UT��y�v#NX�T�4@�\�=a":#/����n��
(�
�Rl��H2/���it�<���nih*�AZӃ�X��sZ�����?ǀ��d��O�b��"@�A���6��c���M~��"&�fW9�u�����J5��v�4���R+�r�� �g�����,�*����-���|a}h��="�w>� ~���{�E��!x���7��Ѕ5ܴܠ����s��8tI��a�����
�ϯ�	Xx�o*���ԛ�W�d�)	�O�b6��g9H?D$6:)��t�mN�M޷�S-y�F�>hAA���WB{�9B	�F��T�B��m�OT��«Vh��W8����-�h�O��c�c�*MK��m�Z���b_��b]�Π� ��g�B��b4fO�1�HQ#��cE�C��q�,�$k2ȉ�G H����a��'���IcaH�NYJ�YG]�K�4ǋ�r_"E��تÎ�j���CZK'�V��Xs�ُ8�o`�Q�A�)�X	��Cc�҆ޛ��*�ՙ/���ܠ������I�Q�!������b6$�kS:3\ceHѠ(���?�MoV �Rsz�xv�����u��<Zj�r���R�������4�n����^����VOC ���aLN{D�>\nC����_iuWp�)}��Q�P�_��׿eV8Jʱ?���q�<�Gh���n�g�$�냧�����A��*`�
���T�`����Sjd�N������ub�ѶIo33���`{�f��I�T�3�Ac
6�&�IݻE�e8x$��޿����:��.H�m��(��l�3}9��=���k�@&�����&n�NWM�qH1���/	��
���ɉ���m��v�'�l�&T��Dj�>KA�3��.4�\���,��!@Xp�x���l�f�*��-M�����Z�E�;I��߹�!2O'ܭ����N뿶S�U���rm�w_��.H�����P�	�6�I��ȽɴD�n�Jc��jM�.�';��p��^����b��CE�Q��h��3��ɵ�j�U�,�[o�ٛ�l��p��m����A`�?��L<׼��ܪ@M6��.������:�.h߉K[�Go[�8�vV2����/�GIu�W��'���PK   �Tj$;�  T  /   images/55269798-4c36-498f-9f6d-2f3e7c8d88bb.jpg�vuPN���.,���,��eqw,N� !���Xp�� �5�%�$������ޭ���qϜ���ꙮSSݏ��� "UEE  ��w��ؘ`R2RRrr�S��A����S�)B�פa�J���������s...�?T��Ł���C�O@ID�������������Y��/7��n(��@�(B�1Љр�h�� *  ���S�0� Lt�?Ai" ���L ��zЉ� ^mLRF>kϐ$��':�'dL6�Wɍ����O�t��fx��/��� 4t �o���_4 ��ш��$�� >m��S��e �_w� �O�@�Р�I�偀��}��=�`��|eAIQ,:�F��3�r��ʍ��L�%��O�φ�_��D��!f9M��J]���>��5Y���TI�b��)�H���:��[����/�T ��e��E|UMO����Vd���_,Ӟ�'��T�������~1?o>��I��t���h�Θ���s��Ɓ�# UB@p�N�BS7D|��?�+u�p���{�te�q�W�n�����z[���N��uN�����d�?��'ax
B�c6b�ڕ���3D�30V�ů[�x*J�:7_7��6ӝl"v���=0�WJ�Ȣ��IF�#�ϋtVSl��f~(ߌf�+����K�Y�ښ�(sP�S�*<�Ό��L�F�|�y�T����T���kz� �]v�$6,:|�*CxRK�~�'e�����uBu)���m��D�Wl�mMPJ�þf�۾�߳�d��T��t�3��3Ó�JK��oD�~� 3��8<a�eoΓ���~��O����W���b���"�/��l��X�䗇��g|f�5I��P1�޺������.M�Q�SJ!�o�j��r�����v���5JuX8����y�6I��2C�tt!��2�:�|ZY2���0�$X@(�D����#�tx�|��:���8�љ�<3-V���؝�ۧ�b>�S�l��0�
�P� �M���xo�f9��zl�z롵�o�d�ld4�FH6�@�K��>۔)���6qP��f�)�Ќ���
@��_+]	)�G���o;\?�
8�P���rG�Ƥ�"y�0^�
?�|"��ʧA"T#u\:󙇡o�����g5ctbi9�;@��͕B�諛t�gr�P�_D�0�����r=���--�<������61��)�n��b|ݬL��e3!���~h�UR�k�m��Sh�6������ +$y:g���=(apQAb>2�ʓH5�9�V�����O��Ι��ΓW��u��Hg�x3�:�S�Bqh��\��U��[{��p�.�o�׷O�g�*B�=���o��:��u=�O{����AP�F���N�ZR��%��7�'؅z�~a�ݍ�s��u���+e#_�DmM)�	5PY�����TtɳV^o(��7u!��<�i6��Ǧ��v�	&��?�,��J�x��+��Z�,$�<�v�����w�=ו�;`%j���٣y��Ӷ�}&��u��y_ݧg[/�]�jn�9�I��L��=�%�#>��t�O��n^��E��}ƥ��*'09S�Kn{eK{\�TsQ��>�W��	�c�@CP^<(�|��)x�(���Kw��-'Z�(��t�f�Dݙ�5R�Qx>55��,s�A6}cU�F.���x�J�|B� 8�4����2)����I�#��=O�-���j�Wԗ5o�k10�������5�5B �Ӑ`��X�gI��t�5�I�P��o����L^p�����:'0
_�*9�xw�h^T�>h�"B���o�=���S���%��G���74�@��T�y�<�3X�a�8�N���%��R��P	஼�{"��U�>Z(����:*�j�Yk�&��g�^6�9zJ�/�x0����ѻ߂5��������t�s�L��J��<qO��}D����jD;�$�{lS��%�Bwa�<����n��:ݚAz��&��A�e4H�ͽS+F�p6�����(tG7g�&\<�^��Ȉ��Gv��������u[�&�sͭ�����£j��3���<_k��ʼO���z"�ƫ8F�U)�NAcxJ�D��j�Q�0OB��� v�Rf[��,k���Y2Ӓ����P�h�1� �)��ɵ|%�@)Zv,(2릲ie�i��&��'���i����y	&�Ԝ�|����-6�{D^	ǜ�����J�څ�Z�b���	�Ry�Q�  `��s�T�}Lg]����$q"yb�ձI1�pۊ�w�(\Z��.W;����r����ag���4��\�)&�aq��^Td��������rsoKՇ��7!ue��̰�ŻXxڔ��� 2Ɇ˯����]�2�	�gƯ������MP�Q�ި)U�N�J70ʄ
�g�F	�PN0��4#Y�l�s�%���Yl|�(i)�!w�y.�V#<�j�����a��v�Y���C7C��F�+��2#Tc��� b��Ti9a�������q2�!�',��x�KEȊ���#��Z���G��y��V��!�G�l������#���M��j{��ͽ�RMeH�	����+Zr�v��u��J�ku�����܁��K&*�ȋ�M��ݞ{��J{�uf��fA�ش{�mt��,�TRF��	����Z*�S¿u����ߴ �`p���"�=�Sr�:��c's��Խ֫v�j<��!����۝�^�j�G����$��V���Ej��F�솛Y��E��ff�)�/i�S+EbW�o׹/E��uv<�<4Sr�N���۬p+k��`�:�A�q|��R��_�Du^��yChrc�w��I%�r$Mz_�]e,"�V0TE\K,KT����1�t܎��dl	aO*���4J&3Ό���}��*���m���^�}o���k~�����HTv=�k;�9\�]�򜵬r��ۇ:leb&����>�`$ 5t�)���FN�*��B*�]���?��չs�Cn;*�z�i�,汊ي��Ee���_g8C�F������Q�s�~´��-Es�WP�PlI�6�
~��2� �d���ٓ�jm��8�^��yGT�P:&����
��䘆��;���_�4��:�zQc������(������ek�آ0$ٻ�@��/�a����;"�p�k K/�3���HRB8���ݦu,�C_�:!:�s������:����ȅ���)K�,������t+E/_P�h�O�ێ�-(�"[I�惨+��W?�;�f� ��g�\�Uӡ�/5:��a�t�R��ln2�����9�>,��{���ڛ�ɘ�ab�>LZzL��DX��[�V�lRQ�-2��&,��Ϻ�$;�Qk41%�j�"�y��^����um�yh�úyB��'�i�6�ޯii�Z��SK��O,�6ɱ]҃�4Q?�j,|r�� N"��9~����L9�� "[?�S�Z�T�� �8!eFʽ`��^�6O�����(��Ȼ�A�ۋ�>�8��Z 35u��_�}4}���E�=�}S�8�b&��;�ܙ���3�r�;���tӇ	��4�� 
E�cv!�$��J�[>�0�>�Up0���P�j1��~@�S'U)�'��廾�'Y�-/@�n�����<(�,�U��dI�VVK���=��ȿ�|%i��A	0�:@M-��1��p�����h��B��pa�n�Y�,��[����w�����s:r=��C�Q�S�*�[ۿ�:B��0�8
3�u=�Ʀ����|��B�6�|n�q�Mݱ'<�7��?��w鯊wDg���v��,���5� ˺�:o��U���l	P�"�pO"|نZkX�P����`2	��B��8FH�2�N�(�L��fD5ױ*M����+���ƣ�'��I}>�P���M-�C�H_G�T���x����p$>qU���9��1]r��J��k���B6��;g���%�]�o>��.����+kzj�ۥ���L�����Oyo/O�����7�����b]E;�eo����u��@б9��DЊ��8�H棭�*)ފN��GΞ1�{M��7/o����V�e~wsv sJG����F%�{V{�J��ʡl73��u��#C��O�oˌTy�>>�ԇb��C�D�z'�#]X���:[M�Y	��i�J]5�/x���+{T�q�='<�	u#7����O�υ/hǤ4����{��i	�BE���x��˅g���v������;�7�J@�I��(�=,?��y�p�,t7��"�����%��?�|5����h�v?(7�ڳ�z��L?bsֆ��F#���c�AduZ_�w�;�ǥx�� �ϧ �9�}�U�'�:�ez�S&w��ך�i7�ו|���oK�0I"^�ﷶ��y)��я�{[��x��Ͼ��5p��YY���ΰ���N3"��	�Y;�+�������'ʤ	Y�1�x�'m(�	g�:���cM�Za��5z6Y��}�a
�Q}q�lv7X�,�xʅLf��o>�+5r++��,�4���yW&��?06UI�Q�a�ٽ8�P<%E��݇p*��u=��w���5��[��G�d�f�e�L5�X���hW"�M��/m�:�ӎ��w���J�ˌK&�+!������ <�E��/�Q˻��,n��/��}��?k��(��I�kX?��Qy��:�%i�w,���(�!�Y|��;��޼�A�a7�3�'�� #�S�1s"~D�1,�>�R����;�`vZ���zR��|���v<�Wch���.��ͪ��z<�E���@pT��	g�h=acU\aE�
8cň�o+�<�C9Z�1�ڙ좩���������B|�w$fX��)?��b׍HGF\"Y�坊/��e�_�;5�U�����z��G�5��sX�ȅ�z�}��.��y���#�|@�ML3i�j���>J���M��D=++n��H���M~yM�-B���)c�e����Ҍ�4��,+�ܝz,n��@N����(_~����x^ 4�U2�
�����}����sܓ�>�틎�4{��N�c��ȧN��l�ސv.I�o�S�u\��@�SY2t��|r�ٞL ��7g26��#��ƒ6�ڶ��6�mr&���#�����
���P��ӂx�xE����D�.�Fk�q�_jd��L�L�=�>�Ѽ�z�zx$`!�p�|B�ߤ�O�)�i-� ÇB'm���)���|��`Q���r�?��\�����#����Ĵ�j�$d�}-���G�L�y1cCP?U�z�LIAܟ\L�l�8&�A�l�y肜��S.��=G!aLPU����\��a~Q	/އ��Fr�Q��jo��=�F:jO�.��&}���g ��x��lV�s�>��Ze��ϐ�q�ʿ:e�5�n�Ȍ�:o6��[:�k���28��{ՠ�3�Z��ӥ%�g�;������һ�V�dAucN�s�ށ��P�E��`Zi*��6]t3!S�Oם�n��=R}��yv� ���KK��P&-`���Q�g^Ʀfے�K�����9�p:��V��%���x?��s+~��_�(�['[ô�V�`}���T9K��`�m�0i1����ّ���ݡ�T�ɳBi!Jz��JZ��� ��%�/�0�"u�#@�з��T�� _��i�Q�Pa~���V�E�|KO:.O:��>3.7�\ȺQ�ݥѴ|��k��9r���/��)2,��L���yq�g����V2�:;?�ʹ�S��oq�"�Ѱ!��j�a�_�e��ܷѰ*�����Q?f����)����@� _=�W4��|S��Bd5��}��tUkf���v��������\i}�f<��q_X����'!z9AO�B�H�d��4��_&H���H���Ϸ��㊥�&��N ���{*��4�j��&�E���o���RW#��4n���PD*��a�R�R�Ky�]��q(O��ЇL��:�7���NJ�_H_c�{Q�EK��(��)u�;�w�W�5�����%�ɓ+p�ʼ�H�L��&�L���?�,��  $�-A�R�WPɭݠ�һ�#>�o��I�~e�2;]�.��f/"ۋ6�1zA��������R����lp[� ��Zқ���O覨_(9��.O��%	�p�پ��]Y�_�����l_L�@+�G��e:�!�퐠�UWNr~��?!S�f�\��յ���B*.o��3�7_<ߦ��Q���V#=�YΈY@ㅋ9���n��x���!wCq�b��%�;��?��.�G�'�"�ӵ9xz��W1�8O 5�Tʞ.�R�l�	�4���IV3���]�ٲ�˴\7��ͮ�z�zT6խ#W��̾w�L#O�k�(.c�O��R�4)��$� u�d�>�D�+s)�f�xE��Pb���D���pH/㿋��oG�{�Ĉ���W�e�k���<K]A��¦�̖�LaiX�z�L�����(�E�9At�vb>%zWw��AT:l�2Z͐�*�|�Y ��7d��>b_IuE�X�I�]ƹ9�埿���xJ�hn&-f��c�]�X�Q	�`ɦ�"I�m�|��3�� �u���yQ����
��a�|���`yib�4�`9J\��b'<�jn�z�}������B��\��KQ����U����Î/J�WEA��qm�v�6�s��eõ�����"'�5o*���{�H����_6Q.��[�OQ�,զ#X��N�7�GZji���}��υ�3�xǫ�w(y���i���<H��Z%b��G ǯ�.��Fښ��`'���x�ȧ�F}�o����}����?��%)�a����)sAzR-��N2֎���%�N�2��z}〔�^M��b���R�&�=s��
Ɛ�8V;-�z8E�f.�	�,�.8���h�	���!��|yle��$o�g��=:��V��?��F�8�C��myn�+_�LB�:v��A$��C�!`��t�H�{]�n�bb��M�A�uh��|R��ťAơ�צ(E-3\��;�}�a{��C��i<��a�!{Dz��S��v�x��;v���ĥ|J�e3t���HH� T"����ٓA�32@CT���B�&�~Vj9�Ko
��I��Bg^.O���F[�Fٻy[��x��lآox�O0�2�W�P�W�C������r_��J0i������>�:�>m<[#!G|Zi�n��m~]R���i�\y�� �����9cHפI~ϻp�7�+Y�.�,����v�H����@�[`\-�N��q�? PK   ��U���[B� B� /   images/b676df13-73e2-41ea-8e8a-dc46dce3d5cb.jpg��X��/�X 8�� �	��'8�aq	��]	.!�]�-�!�.�.�Cp�K��������9w�{�ƺ~S]U���4��
�����    �xZ |�|���������� ���+l�W888�H��HiȨHIX_S��SPr�Y��оCx�� 6&&66&.6%&-!161&..1.>)�KRL4ZJJ\,L"\B:"��� <4$�$Z "�S��#
�_��{C@DBy�������^A~�4�DB  �"�>������;U�-��Q�)S��o]K�r�ǂiD������aR��{�b�3�%�
۶�=֎�nbva\,�Ԣ���;~/�*����Cp��9șɖ�+��?z�z�q����E��8�Y��
OA��Zc�P $����c9��0�/��>R��h�������ȡ�$�w:-�Z�|sv&��|�]�y0Gd��1!�%&Q|�t{�KmA\�<:����b��� sH��o"�ϟ /.A��C�B�)���&���]�D�DźD�*�im^���l���z��ZMS�Q���V̓���ܼ`�w�U�{خMaĴ��p�����`|{�6.U�L�T>���Ţ'o#/�����*�fİ�����`�	O��X{�n���GYƧ���u�	�:_-?J�'^����jo�l
�Ln
H�/	�OjhY����v^��G���k:;��3��9��J��cQk	��FQSF�mI���m�"��>/&��?�1�@$�����\���Z����	)��^õV
L�)�CU�!����*'J�# -Z��LV���6�z�"����>p�.��HO���BԂ�c��rH�zL��>�N3��!����F�ي�ن�3��[���P��k�T�;`�s⯇mF*;	�"�^��9H`*5���	e� x�n���EN��"�t m���G'�3ݯ#��QGQ����Q!����rxٴ=�N�[�۹���2qw8��X-@I^�IY�Zh�&�����Tu��ǿv��N��d�d���Oj����H! ��$	�X �y����
ǵx^ċ2*3�n>FmW�g�WP������4Ȅ"	T�j(��_m��hn�(��c�L�d��0����]�k�05}g=��*�sT��TҸVXUM�P
W��7":��	�����4)�t!����(J�>�珘��!�O������А�)mzO��-�����i</	�CD�=�b��,\0�C��b�2c*q�C��a�av3��9��s��`4En���"��	iP����ͽpEH�InJ8(��ө��@�s��y����1Y?�
6�lBbdx�,ōȐ�&\�>�׬��'��q��ݳ�F�m���Չ�x�!|	^|	�e9�}���{&F����%�hȂC�]�_�4L?0��! aq��vx�ΤqϞ�GZK^�z�}��dB̖z���+,�u~������Sӳ���A��3�Y籃}�^,�;'�h��Qh4��py�TF~��'�_tN�^�hړ˳�L��s��V�ujm���FϠ��$�����i
X�����1��x�Y.����Z8��$�k�?4�l����뚽b3����o|�]�h(�ĭ�
�����e����(�<����}_%)<䀖#L�TK+�8�O3:h�l���@�a\��K�7l�F�lS����$�mN���కڀo��4��Ӆ���
P@6y�C�&?%X��,5$�S��P��N�G�
N���Z15�,�����y�+�-�Ps�u$�g,^3���H�P��1Ʀ<�k��跥Yɱ������L�u.�J<�4�Pg�^�'�Ha��6x�PN�Z:����j�M���6,� �06В��e� �<5-��#���ds�u/�M�KK�	��.��i�0���2v_��;�+�e��L�s��{_�^��;��������Ջ��M{BE�.9����3x�KR��_5/����H[I��d����ߠ3�������>�[hx�OG�,�}����U��m�H~��d3b�<*9�E����tg5��K���Y��n��z�{�Y�ŕ>�'��М�7��+������y�ۖ�~�4����kj�(~?'%��ng�^RY�vL�x���x��ш���=	�� �i��=�D#H�%R/c+e�؀>�RLI]�D�߶���W��W�����ޏ�J��x��W11��9�cC�)���\�BU8;��v����5�,HfIg��{����j����N��֣������F���h.mn)��<�[5M�N�N��H��K��'=��Jb#zH	])7�^�<��V���217�4��9�n��4���Gf���^J�ĢP����b��d-�QK&|,��H	q��^�x�@���Q���{V�����NQ�!�̒�#w�Z�m�D��x������Ǆ2>��H��&�'�B$@����{��)����J 46[��;�AO��[���[�89TB�4_w^�ȑ���ZY`�.�ҿ����2T�_�����F�|م�4-�BR�p2�m5>�7��T��z�[�X��v��.�%Ԏ���Z}�'���ʂby�;\�A/>�^O~gj�T5�����r�Y1��z�jz�J�C�
�>�j���L_F�����v�	�Ra�!�&8���oY�Z�t�����>4�t\vy,m	q͗qX����S���U��h��bP%�����?&>�b�Z2{cd�<~�n��ʼ�)̑ϸ�-��0�_�*��S�"��=7|�i�����wR���.���̸C���q7#�H���Ğ�M�m���p;�����cEЃ<@�:�^����aV (TN��9`ة`��KBۧ���k��N�����1kSLU 캩���k7�H�b^e��jg���ϴ�9��Z &^���|�9���ʶ�i+(_��J�Lt�yFy3^ˈo��)�h�ܚ��Ȅ�[M���[C.s�K�ߝ������	��?������^7{��y^�{�gL�i�H��p�LИ����ק�P�L��l:g:����ͫ�d������\&T\��d)�ڃ�WarYܔ���߉qL�ڳ#�'�V�3�H��j���=\���]�|����2A�L��O�Rw����_�6f��=~�71�ޡUʙ�8�]�g����J���L���]�����=.���߱�1��{�4|�	5��爰Z2��RU5_m`��k;��xH}�)���)vnD&T=�N+P�T�alRm����n3����,%#P ���-��A/^WP0����6�m!�-�-\�Ռ$���>$&��Z���ߨ�!�t��b��gء��x�8�X�s��1�3q�(��aؼ�p�X1����*����A�[ͨ�$��ʹ-��/��*9�ך4�8��V�=��z���>�<����C�k�Ou�/Gn$�3!<pC:JwC!3c롵�?h�<3�38y#���
ɰ7v=��-U�BsU���^���ڑj�&k���`6�r���\�]�tJ��-FO������W�(ϯ٣�Z�<n���lD��s�-lz@Y}�O��Z܅��5��oT+�3��h7���}��~�I9jx�2�L%�Qp��^�m;�S,͓�i����F�<��*��c��s���7כ\��Y��ÊO_
�����.��#��/��_�m7';lc#>�ڿv���qQi�Ҟ&Y|��rq�M���/ﯝ�b/�;��Ԑ\IʗhhxH7��Jk-�ڭ���`R�w)���@���M�e,�	/�5u�al�Y߳X���	��gΛ�=���eݽ�Qz��T�	 �<���Xp�s,�Ρ������>tu:�r�OT�d�v��y��)}Ψ�U#%}�5:�1�n>����g�\n����}=ɹ>��7�ܖ3d.���(���9�x��s`�q�A��q���k=��)6J.��*�h2w<y�F�	�MW���9��~���@��V�VK�!�t�P�o�Ls��~B��ּ���sx7d�o깛��`��(v0�n��,�T�������Yϣ�_;gd�����~6Bߋ��'�<q���t4�v�UЮ�s�~B�N�W1��pGI���'sJ���g���i�Ø���@����?[��	��s��'���Hz��#v�g�����M)(K�Ԭ���J,妉�&tZǐT�|_D8�¯���]�Ӹ�S�
��߈�eʙ>f�?rIj��v��:�֚_4�\ �ᥫ����{�������k���I��hY�tU���9mm��=�S?Z7�ehh��y����/|Y)�S���cZ8�RW�N��[E3W����$n�t��gR?�z��7�To�~gx��VL��B6G"Ķ�z��Z�k-�wE0Ýo��sXS�Q��b�Rbv���7�D����r��)�J�
��cRp�R�����$����E���m�2��/&����O#1�y]��0ãQ�:ļ�(�|��)P�f1%��!�����29#зs�P�����
�E!CcS�B�L��HMgp��7�`{��#	Tm�|{��}\�i��]�۵��-��9�F*iGSO��O��a@���L˧%�8]�5�~q9��y�!����k]�Ny;p���ތ�έ e"�(8Bm��+@���h�Ӯ\�ׅw�:^A7+ 1ʃ� Y�t���O�gx9B0�׃�3�,�{��!�B�KB{�3�Q���z��~ǲ5���^��hw����\)��ʃx�0"&��-Blb\mR�ވ!#��V��s#r���~�R?�b�5��u����%����ȃ�<����YȂ*C�U%P���Q�$e�Ij�Ë���?N�Ѭ�}h���Ռ��H^�@�՝f̬�Ê�eC���_fnǂ��K�j�rd{�vf}pD�ɽ�ZG���g�o��nD���S6{����v�ӄ'���u��k�o�q$�VRiЙ��Gq)�(J�g�hk��i��i�^�Ɇ �:��;�g�v�N�!F�F�l�����K��>vD��y�K�ڥ�D�\�[�h@! ۳�۾���4��vޘ?�1�o�#�L��Y1b-)�n�����,�^��H;���N$�v�<v3�.k?p	"1	��BYx~���f���`��J�"��H�� 2	�T���|�k?����R����Y��	���O`GCWg	+s��_�`�[=��w�vБ6�sH�M�N��l��HhPq?�8tNi<��`�iρ3!�?M���|xs$�i����f�� �$D&�CG疤(U-C�BvBeS�◢�N��(��gL�aBg��u�Kg�����=���P��:?>��ۭ����gj��M��sk����h�J����o=��U�7̟ ��AE�px`x`NtT���:8��R�XC���*��!@�A�N��� Gy!�ܿ� �����K��G�K�Ã̢�5.�cD%ҌftN�����w���<�ߙ�~IVJ�/��|����S���l\D/�Q�i�&Ӡ�d�ic� J	�	��gsBKQAY������$Y����FF�5lӄ�9�i(gd:^�qbq��0�$?�s��W�܅�ypb��ܽ�2�:*��	Ѝ�1�������p)u;.��kU??��Y�vH�Ơ�i�9�ʄŪ��Ƈ��w"���v��h�:�;��TD3����`�߈��Њ��YX!�Ԧr�1�i���S�DV�cq�5֧Aђ"}����n�zN��Jc
��X�ц�� V�.[$5�Qk�Ş�:�C�A���gAg��L�e���r��x��˙ߎ����'����D�r|YJ�h�V.�}��r�r���x���Q��+�,�ё�}jح�@�[��В;��C���n�^l�0a7��*j$j��@7�$5�<����K��x�g\��.z���]���{	{݁�㬛�B\�W�eI&
w��)������[�Xٌ�cJC���I�e���i�J�"e����z-{�z�p�ޱt�^�7�
/98��x��ѽ8�0aJ�-i�5)�]eie~�����VoGZ�9�YoF���s=�7��:���a��aL�$�N�	���<�5 ��𺽉L�N��}?9os�ZA�%TTO����9�\A=3�R�6�)D?�a������ӷT�N?��D�r藓��`�<�M�F6�&n�G�<O���RA�(��?���in͟1hk��[؈�*�ç�*X��8��V��fU�~ts�LLoQG�I'�W�;g�9�B����2w�r覣Kc� �؞5Z��Qo�4�:�7�7�5�BuPT"�H��k2<�ϤL𣏕͞'��4N<p'j�>X5�kl���הʧ,4J-B�?����ZmA쉴�%�ZZ���\ �2~�Jq}%�1&Q�^x���#J���u+�
4�c��Vs?͞~�9���jYŞZ}ߑf�ɗ���B" W5k�$�G�0���W�Y�@����Y\�,�����ꠝ�^�λf��osyt��I�H�V�~}��M`���~c�����
B�W�h�b�Wio�����F�2��J[=�v�SQCn�a<>�w�/��=.oM@�t�e�!Y�����|�H�E3�����t��f�Y-S�R�]�����IkPJ{v#ZN-�����YNz2��K����P�DK�g*�,t�����Ev�����ԪC�3�_��Q"��3f4��a�ڝp�q0ngT�L�m:u2f�g�-Yr �WLj�m�YQ�^�ˑ`������Ys��#;E��2������T����,����mD�@x	�[j�`�!a�!��/>��n�ǜ�4�R�ڴ=���{�(��������H8�x�r�T��N+�NՒ�k�=���B�����؜�'���n�
q��!��D\i�*��_C�|:�@+R��4�+q���"��M����:2�6|""p|��BJ�1t��Y�*B��9���&���ˈ�� ��z�[�Tι���gu�[��EL%V�%y� �CC���H_�7%�yGYl{��eWY�,�{�i��ɣ�l2h ���ߴ���̢���X�k��B�_z
o��,�.b��t����]����<�	�,/�驺W&��X�1����,l��$�Q(���J��:$��k�c�ͣ�`mS�
J%;�ސ�BM�e4�E���b�K����0�29?J19���E�(TITL@fV�t�g�A=uI����t(άy��BPF�v�k������T�R�����
`
 f� ³h� Y���sE:&[@֟؆ْ��y���i�R5�*�^�za/KBҊ)�s�rV{��rp.vVs�&��+�y����XЈ�4H����m���?א��H*��h*/�C�7���ܐ4Ɵ��1v:�_�{V݊y6���w����_�??�����<&1�5Fp���m�����}uP�D^���&�$��h�����*��L4K�֥їO�+� �v�U��M�O Gk���&�c.C��ƀCI���B������OV�ӱ���@p��A���?/ ?ϟ S'7�s;��|Q��"��O�;���UC�C���o?�0�$5��φ�D6<!G^��wt��CC�:�^���r��^��Q��Q5*�e�Gs+#�mL���{���� ��ڊ�'�{�n6��'	��H
n~k�Ɗ�'�����=tU�z<��Ү�S���@FFADA � � $d�W�q�9�hh��	ޣЉ�:rK��ӫ|#i��4@Cx��	�	��l*!��C[�%���C���+�2�NX�T}��Li=Hݸ����\��N�.,H��1����쿧�7��e|��~� �V���k����=�A�>��@�<��_�2�!��NF�+������"!�[
�jЇ
�2�l���Iw�!���2����xu�n�r�h���GG�[�'�=�l��x>��^��X�-נ�	|qH�Һ����+�]�Dp]�X�����,��_r���F��yl{��b����M��RnX����ʼ�JV��S���Jv���<�k�t|<ޞh��O�DP�l�f��V�)���pg�^���Λ�	��eN4�G�A�"W;�}�r��-^F�8���Z��5���V��9�m��FɄ<�qM��z��K���ޣɁ�Q�s*o}:����y�F�9� ��*
~,w�-�ms��	�1)$!�g�o�q�X1������	KAӂm{�e��բL��G	��z����6�m_I�P����(j�;�J6�]��`�W��{&�Pta�yR�F�JP͈-0]a[4�䊟.�=:W���|Dr�.�;aϥ�
�����k�����%y;�8���#xG�Z?"x5=?-�8��p��V[��'�Q�O�� ٟ��li�Lp{�Q?�B�Rk�����',�X��U"		���F��A:y.ljY�lZ�ٕ���Y�C�������$���4-u�����I��ͩ��8��b]�0�m�1�#,(Gޯ-��zI�:��5��D�b�Q�r�
�=�U�$�bM�᤹�C��N2��)dCl�ʊ�槻@T?��j��������nD���{܄�DL���=��_ݹ��k���`��g--���2��zK#�#��(UN�f���j_{D �+A\��IR�!l�h�e>�Տ�X����'���@c0�0�O��R�W=_��zo��g���g����_�k��[y�H?�� N͢IS��?��hN��bOC�8)G=�B:�㦗��'���^�v�
�K��7;��E;�EJY8@Ck�/|��ً�n��bG�PO^�&i�}��,��)�����[ZX�@7���a��}b�3���B#���HD����m��+yu�W��Z	�D
z���&��%��Z�ߛ�~y@���v^?���v��3ö�cpHz�_��Z+�5��q�*��V����&�$T��lc�腉5Ặ�l�@��Z�o^�-ơ�����Oa�|/�U�l�"_ǂ�'uL�/u��O�{o2{�4j^e�}7���	 qo*]"�A@�������H�a���s���5`;8縌�j�̧gI�����ƿ�h�;Hj��-W��vy��7uǥ�����Q߬ғ/�F��	��Y�1:$o��I:ȉ֬ٝ�mq�z��o�ZI�5�7M�&�?�5�E�UV���;�cH�=Qx3�g�Š�	�	C���[����M�@�ӫ�h�7��d+ә&�:�["�kM�%�Q�g�� ��"e��~<Y(�?��������?c�o{���p�;�%��4rN�9=�cR�wt>:���%�/#�~��y���s\���TzpIq�@<ԅ3�*�/�`[�(��.�+�5A^ڽ�d�q�6�	%��BJI�
��Rc$��<��$�`�Rb~id���G�Á��^��j�'`} 36b}��0ݯ�I����@��轁L��I�)<f0�_F,��`E�οK<-Y���1����Q�vdQ�|]U4u���pU���ܯ3�L�6��|��+����H���Xg�\����c��҅�6��)7X�Tեv�Ii�X��gk
����c��/��L���bK�9�Ʈo�	-��8����f��%x��ئ"��'R,��� �Zp������>D�����P.�^Nb���ABM���yZ!���
2��V�h6���Z�رJ���IM^�\��v���jWv�)��ީ�8�T��w&hJ�e^/�=�M�z�!6l�����iK�W�?�R�`�gP�� ,��v����4�6�Mֻ��{�.�CB��a��
%��ͷn�j�9R*>�w�|�����o^Lq��*w/2:7��X��c��"��f��̱���]
r�R��|՘�{Uf�����Z?$�*�Y�`�R	=��B�K:��j
Id��i_�Je�T#�f�V�x���S�}�����D��!j�k���,ѺS&hi�&���V������೨�����,����I��AzFE���26������x&v:k��oӭR��%;��j1�����b��L��U\��M�*�����XJ4[��� _F��m���ڛX`FáƔ��QA�2�*���1��knS}9���j�.�Q���4R>��3'*3�Q"�B������"�	f\-?�#K�1���+]��æ=�tw� j_Jb3g�Sz��)��O
)L�����*@gٶȐ/�{{i�s�9��K�S�gQ���r�3=�w#����:�Lhz/&"�g��=�C����E�!�� �XAO�HSZ������r.f҈�k�/��*��{�0��B�����SIߥUY��]]�1ȴ�ZF�	�U.]�
�4�����Q��oK���<�s^.'�+fE�˺s� ����R�jh�.����,6�d��4◟?��%~�6�)���@
��Mr��	�
�����ӫ	V�a��]��W�*93tN������V�:���k���]KV������Ӣ�mA�{���fi�k��nxF]L��h����n+��I=1�~Xy��m�n5���[�b=��7n�@��>��h�}tīל�֭�]�bX&�C4SE3R�;�o�6�X~G�z�q��k6~���9�
�mAQ<�i�@USWyk�Ѕ���Kh�� [ �D�J~��]��l�d�X��8�̷���z�rF�ON}��O7�T�H���z������őeci�t[u�9�eN���q��������x�8Þ�O>�pK1�W�!q���=H�(`��k��K���׵���J�}��B<�?�;���`��@�ϡ��������u�i*ZA��H'�l[1!lϩ��Xڎ^r�.�:�yWi�?�-Y{�y�%Y[�V���Q���G,� n��W'�p�k�����0����Z�[�1�߆wȹ��dwf'�wOe�7�UQ�(��R�&���2/�%N�Sz�Ǯ��2oNq���Bәp�Lᔬ���7�s}I+]ջ��Ǻ5/����U�A ���s�,�^O ��-5��[V}*�J�dq�o����d�%�k�N�\oG�L�hC츐��?h�
X<�-�TV��El��M����Z������}�;[*Qd�U�Z�=��q��+S	_���*�"��ɶ�Is��3vXԍ	�^��؁�/�Q��}�De�u��g-��Mz��
���h��UӢ\�V�����߳����2 ���%�Za�׽�D ���q��E�2D�%I���^g����mΨ�<��y� ���{g��Z �;G;H���V�v�3�l�ĴT�~��`�س�ƪ�|���AG5�zEN.vPM6�'�cȽ�ye��-��↷m��_�!���_R[��ɑ�`ty»grѪ*��C�>�a����Y������+�נ�q�aA��l�u�e�`;e�����4"� ���D��^-,��
U3i���gF}�l �7z���,A��u�Xb���8��G=��E'�}�M��w*%���4d5��J�p����r���J�r��݄��Y ù��)����v��{��259N�O�Ū�T�����1���cZ�ZT��F���ܹ-�Pg�"���x,��&^�m���~1��=�I�d�̚⫄�-$Ai���46�b]�,�g5��g���s��+Є����3��3D�/9��uG/��8��V^=9A��'kfZT")A[��ĬOZ�oj�+vx/��Z�孎$lj�E�Yy�Tز�L�J�?�>���R�o��3����ix��L y>6���)~�=�Y'�B��p���D�\J6Q���'��}��>�����HA�ՙ�1�k��	ll2�FBMk6ַ{�:
�D?3X燰�	wC�?��.d-�r+lC-"���?��)�խ�V�Q;#27�Y4�b�D-�e���&}�v�J>��P��kОX	Ǥ\mZ�-�E�TO���U3	)���W�y�}��^-��l�v��w�'�?&�.5���'�2�@4��)Q��8�N%͊g0k�M�Ѩ���P:3�X��E�<ȐR�QG/o��sE�������!��!)=�z��b"Ӗ�TW:gAM��Tk!�� ^)���R�ћT�O4m"�d���&b��v_MZ`,�_����Rs ����9�xj�U�;z<2�i���<�{y��	-�(ZdH�iG
KM
qD=�ص���8#t.D����:\��<\��?���LAmD�;eSz8w�aZ)O����K�$WQ�'����ߜ�8�o($���T����Ŵ.OJKm�@ag�w&���@kM�*D������#	ς��6^�up���r=��V⋇U��`��fpv8T�b�9��]t�Qfא�QT�ԗ��*�����̄��.���P)a�bn��G��A�sN���m�մpsS��M��ߡP�_H����Ɖ�� �O] Xc��K,Ja|)jg�J�m$qUz6�`򃖦�E��h���&{��h��l,>aMY��\�4�	L�8ۤ��_���&�`sB�����Z�z��@0�<<V��G����n���o�j�W����m�X�Ŀ���)�\N[ɇzs�-�Y��~�/����h:��2��f\X]���g3j@������ʲ4|��'�#B�G�:�1�'ehڼ>5������3� i!��� v��^i�^�߻�TC	�`C�6q��`�u�/�Csm��祗��"���z�֡G���mѷa��:��  ��l&-��k|��ؔ�䎝ZyoY��M��������#CcN,�t+V����A	S޾�^�ÚvK`ڒ�,(�g%LpU�
o&g�_t�Q�`x)�5\w<$ZT{76z�RF��B#Rd�ޢ�'O��G3.P�\��䀨ƭl�L�0�XW(��Ë
��A-[zD�w��DX��K����_�hZ�4��
Q��e�u7��
�c?rQ�d�V��@�|�^�[17�ơ|�'�^Yj��4vө����m,fe Z/���]F�`��l}4���3Vq�S�r�v(-�>�����94~1~KJ���ٯ@�6Pn-Л�sN�*#q1z����5��q��$]�={S�g������:���! ·�JL�I4Y���W:�[��7��N�4�=��n
�~ (誻���\�C/|�[u��t����M]Ή�W��I�/��4���G��]5R����8�ob��6��ci��l7݇����od��"|�9@�1sy��! �!��r�	O��ޟ*�;l���#	�s�4SJ�qg�=�q�d�TF\�B�[O:�úD���ٹ�*R�f0Hj�rq� �l,.�0�r`�g��![����,�ălR�w'C�����E����*��%Ry��ˏ�NG ��y�	�f��� d��eL�э2->͋�?�;)�A:�5 �K0y��ß���=����#��B`[Jn��!N��pivs-Cy��9#�sN��'�e��3�Vɔ�Da�l?�g�ÿh������r�(;o#��M��T��_ ��@���ߴy�!�i
���=��HE[�f^â�q�&�)���y��},����|\���a��f�o��Բ�|v.����dE|����h��/�37ki��p!��:p�#ё�K�T�?���ļ
W�l=���E_�Yf����&����R� 6� :�zabˈ���@�Q��C�rKZ���CmS���0�Z}DW��7űS�G��Nȕr�W��� �%��v���%�8t�x��!���R�\�N���#�M>CbS���@	kQ*˸ys�g�"��X�XF|~�y��á���>d3�x�w1��[�O��8o�_B/��Ɲ�)����M>�C-P��B��Re�bl��5~��l��|�s:|��Yy�s&�dd�bS#v7���k^㟛�vd�ݝ�&��W���t8b�5\.�j|k#�ۂYs:��.08%X�I��_����Ml܄pm�>�Sok����:�ِ��#^Α�v�'@!\�5�6�L��	Pk�G|`�~R7���%�ٔ�Z�@B �ܷ�K�X��_X�B��v���I�0�@����d��A��<���䙨�g+m�8��Kߏ���^��ф9��k[ڽ z������/�t��9;L}@l�Q!���n��sV�dw����C��yt�h�4���D�ym^�RH�[�X�[k�	!/bUD3�c�O�ݲD�bB��`��H��{�%yo�L����}�6������2/�����`K���9{7�^ ]ш��­�!W���Uyv�Ne�aƭC��T� �����H����O_g�fu�.�h<$��-ڴ������ܫ\��;�]��..�Z5*-[��m��i�E�1�&��d`L�{o쐪_��� olT�>e�� ��t���G��^���R���j�i�ښt����f�ȮG�8�b����͘I��<�
�pT�D��G�l'f�jVݹ����|�E>�N��>�p���^y�Z�������(���%�"\[�Cn�L�a��<��n�ئ����C����S/$_�\e������Q!_�`���zC�0�gv��������P���gT3�a)\�bVqh+3��*=��P��n���&p�����i#ul$Ax)�K���,��8Up��i�D��2@*�t�W�%L8�<H�iJi��6|��y{`��bWnH��v�ʘ�kn�l��Ԑp^`F&�=˭�g��U�����tJ=�b�gA�)c������4��i�v�p�*su��.ٞ�Maлf�R�rMJ�
��m�ѳc�T�I��+�R>ѵ�:��\b��yT�׌��"���p�e����$�,=��b�^.�Fd�� =��9*�<����+�n0U���:e�kN^��������F�&���-����xm�I��4��[�.�#l1.G�*q�N�INyi�v	պ��H�k �< �@�[��*>9��$R`¸W�CZ%A�-8_d혁���~Bs؍aA`�9z�j�5�y"�I�b"+�_���޸��W�Һ$��Ե��H�9)T�	r�~uݚ����ǌS��?g{e�(�+���l9];��U��Z���Aԡ������ݺ�of��x�����*=z��y���[؏�[(����(��՛��>]���{�9}H60x��e�	$�F8��-�.d�an�L�6�2k�
�d���1�c����|If���j���3K=z��tݮ�*Y��Bf 	 �re�M�%XF(�i���Zb����$��]���نL���%@}"�z�}1�<��i�D�R�P���k�+��u,~1ʀ5+��Ջ!R`��{�]惿��H����������d�E����,��C�>��o�w݆`��Dc�������O��>�N��}��)�;���~QY��+3i�+��0��m~]��svs7i��7�'ױ'�xY�f{�=R��]J>;9�rl^��Ns�'�7w��\�N�1+��L,�� v-X�z�{e�|�p@Oh��R�����s���ra$��\1�=1ֵPZ�Y�&��}-p�^�Le�k8_b0��L�U�幆�^��i�)��NS��{yץ�b;'鞞��dB~�O!LL�8�>R=l6;���C9���Þ�E�j|�pŘn3ۭ6�B ��F��A����퓳?6�������{]� גM��r/��?<gq2������ZT�}��Dea�^3�>[i���$_�[}�Aj���E�h�Ǡ{Q(�C~�9���	��LO)�yd����Bv�W�jf-e=|�����?L�c$���o������;��v�V ��G���&\m?6Z���o{�h�0z{=%u#��N�q��	�h�yf�Iw�K|�kH�JQ�<-�79,��K���T�-0�3Dl?���]�E�OW��j��<?'�*�=�j]EK���j�a���_�#釮���5(�S����S���j�i�J�0���q�!������%��t��9m�8z`��Έ�$ø���E�
���ݲ�T�����Y�������SR�,S��'x�JE��������y��y����@�ԡ��3���|[ �39u�(��#ӻ�/火��W���n�uɶنqU�艱�iUt(�G!�#A+9�ѺJ*�b8=�Y#��#��J��#
����*a}ia�i� ��wFZ'z%ٴ��8F�z%���E%�h0���%y�]@�[��d�����q�d@X�C��(��S�dQ�	��톦s޽^���R���2������Z ��L<z ���D����g�]�������D��	�	���KϤ�LJ��m���ڿ���' ���B�g��V����'�g�רF/�9wo|:�8v'�e�6��LȈ�7_�P����n-�� q��'�[&+�����GW�$��[u��]m�kޜᯜ��5��?aY3o�������q�OP�Z�F�7���������&)�:;_�L��Ѕ��󿄑gA�_�����?HN#��y/�@�Q�RD���篖�k��D���wD���tt���̓�f��d��������o��E`�Ү3HDT��?۽EH�ӄ����2�q#�k��X{�8c�mxqww�Bqw-��E����k���C�Rܭh�������O����w�K��s��=I699W��f�)ϵ�+f�D��������x.1sE����U���hW"��C��x~"����{���5��J00��ٖ�g�՟��C�v�����}������tT�A��ޖ���,��$���%]���MMձ>��ڲ��!�Ne۽n��Q^t��2^#��7@Y�/Gs��Ԧ���M3��vۊ�D|��(}7M@mX�qtty��0���#�O_���Tq0 �i�х\Մэ��!�x�q�Y/v�fl�@� ���R$Ց�\lIEyr$��A�����%OhyRV��hl�:�&��K����y��e��ѳ�(�Oe�خ��θ��z�[v� �w���~=S�z	�LM8{�2|�=$^_g$��!B����(|�=W���RM�k��-le�Ê�A�(�q���|7Q�ny�>�+����u����5#��=F�w�-[��b���H/2�bJ{ޗX����K�*�Cڡ�����Q���|�/hz��m�c��9�;N�i|�$�fVG�] ���{R1/ꉚY�D�P�)1Ŵ�ȰE���/`Z�c5����ƐL��aҺ�n�3	�@�
KC�W]��=�b�2?s�����w��g�����P8ǃ�F[e�{�8[M�g<o�����Ħ�ʞ���Ji����*�����2Kx.�F�İn�nlyH�v�Érպ$����������#���ZX�wD'��f{~9v�*,�����%x5��<o�i'#��B��	 ��0�f��5Z��� y��{PI/�Ukv#�'�*���;���WXoPi����<�
�&�9�+���~����=�s�?,ǤS(>%��$�}+���wjHC��gw_d+�s�4_=b[A[�Y)�i���2�n�g�m*Ջ�yڭ#wt�t�m�B7�JQyq��4�:~�!
�leOc@<�<7�2Ƶ'�ӄ֖QpQ˸Ņ��V���3��P�Zv=�XW�I�x����5��,f�/��^F����֧�0�-\�_D'PL�/��f��m�Ip�vP���?:WBEM���W��.�.��7�f�J��W�#{*�^�J������^��#�E�p��ٍ��6��߲��l����f�����:M�w��?�j�!HP`��n�y	�N�]�Ϧ���}ל���ڵ��Y<�9"���S�	$�'�UO0u��!�a��_Oۤ�����S5�f��������]�c��0`Y?���<�Go��Y�܌�멲Rg��h�������ʨ+��?�6\�|DN���'��̰���z�+�@g�('g0�LC^^a�e�ɓm���[X��l���|YD����:��AU�&S��j��1��-u���w�������FJ��b�P�����vs]�WgbȐq�����[LrF�g�aC�p�T�r�rsk&�rj����� ���I�.�ќ Ņ��k��et��!'��-�=��{��'��;3��_�'��wҧ}��DI��]������;��F��|c���9v���Gz���4�o?��8�;�eM��t��͵,��O{J{�gK%M��K9���i�����B���C���I���$�eg�r��ú�����Q��da}(�E�х��R�TYt����h��S�OA$bb2�\2Ώ}@�P��͛zp��F��c�|�3�ט��H)�4^��
�o��k���'��y����^b�=��Z�r`]���h�]�(��8wpɑ�|ߋ�d�� o�CZ�麟!��ڇl��>��I��vb�	؍�+4^��Ͽ���h����{�}��?��%7����ϊ�la05��>!y<YKڄS�2�Ma?Ǟ�~�~���ɖp�M�!W|�����<q4^x��ޘI*SlvX��[��K(sE"6��+<v�2Uگ���H�R������ �P�p0���0�u�ֿ��X�8T�⪰��� �@\I#��
���B��%�
>�zL�EӢ]a���@��b;�+�Ŝr����]G��C��E	=3��rk�~�z����Ϣ����hR�o[)��H�n�I�OǊx��
��^�sg?��?����jw��s�C��5�T��<)q;!�oЂ����7gW��d�4��b�� 2C��2��O���$�'p��iY�i�ww0�&	QvvD06Ќ��}{F�<��z�n��v��s_�{���>3�+��b�=� T�?��#��&�H#t���p ���=8e���܈��8;��"Q���G��P��\�7� �1 ��n�{v��f�����9�������� d�OD��Hcn؀��&;�Y;s�fK<��q������9%Py�3�}���E?����h�(���z�1Amή����՛NU<���+�u��⠊�����Oʱ c��f���u�c^߮X��[���K4.��˨B�A�m�H*8d6�ɷ�:d�ź��V����ص��W��>#�J��J���
�>�E��sx:��/�b����ܱZ���Y����`@�����d��a.$��G�'k1��B
�2�K�����������
��w�d�����
����]���N8\Jv.qLjNUZ	�@I�(�?}hD<�>��z��ͣQ��h4�� ��o��q
�e]��U��l��;iܦ��;��Nga2�=Wh�$�6i�Tϋ�R�Ww(�͠N������K�]��5Rʢ�ۮP/4w��_����CL�z@�6:��%?�=�lo���W�Qi�M	��݂s�1K�a�(R@Q�#���aq��ǯu$����?��=-��LΛ�Ed��w|���9�.95a��tY�PF¨��~Yxw^JFJ�RN��B]!��=GZ����f�ަ�U�I�����K��,9iߺ��S>٤ƈ9�T�|Ң��ִ'�ن4bV&����vgMr��t�4��q"݋\$���?�,���w�L����?f9����.��9}�v����ڴK�}�Lk��)�Z@��M	F؜�yCk!�?YȆ!]AԌ��˙����2�p���w����)�I����z��� �q���'��ߵ:e���r.�QK'G���"EJUɷ��Cղ��T�o&3���9KS8v{y�+����e�������T/2��eM��F��v~�<�9���״X���&hBoI�(�n�O]��n���CTU�=#x�L��FPEȊ��>m�K�yiEXR�s-�[Kƞ���΂?�5Kua\�P{8���T����3�`�Ї�pH.K8Y�����^�~�ǎ6��m���+���vB7�Jmŉ$^�ŀ��З�wP�H��7��It�	جTԇ���u�%Q�a�i_�v]?K�R���$nMTP��&����+����mS�������	�&�h�E�H5����e��o ���y��0�[�8�婾>�Qi8JE�.���GU��X��B��"�.��!��� 5ӛ���O=�[V�u��k�r���U��� �(̯zKGY".5�7�m��y����7�QDn���g�҈�#�f��-i�!^����P�_�NMH���tᑋ_ݢ���W�̻����o#d���<q����ry����G$Ԣ+9G�15����]��~�����6�ff#L����<|�:�(�Y�ku��?����񳣩i�X�;	���z�U�Q�w��	���@�����������~Lh,�w>aS�����SP�dA}�湸s0��q��aa�l���	�K��V���I�y��@�-���
_IJ�{�t���$�j�p�%������goI*_�\��qp*�3DdE]�$#���~@�����Q��FkD1@B$�o�P��Y�O,�0�5�l�4bq���`'$�5�Pg��?�L8������{$�S��iD�ve/sЯlsc�M_�Ͳ*��Ԗ`�e�l���eK�x؈cn��cf�@�gvd��H����3a�6:�.i[#;��b�y^�,��}n!��z����J����]sB.��o U#{��*��
���/x������;8(ae�_\'$J�M�U�?
�Wk͘�v*�2�Z�,Ř�� ���Z���`�)A�������Z���S��y�IÖB�6%�gY�Ѹ��A5�{��6�5zn�#R<u-n<��V�ߕ�w���|f�b��lb|ܔ���WF;����q^J�:�Ί��B��2��٢N���x��VB6[���BgS�h�R����u�߷�rG$� s�mQ�+s��b��WXx���%���\1��A6��2�����+��	�NUV�"﭂�P�����9۬5H�yBǼ[mϷB��M�u���+�[�&��k��\�^O���W����Z��.l�����7���g9��x�N�ǖ���vp��ǵ�5�j!Ge��qZD�h}�Bq��4���o���6L�
���Ř�N�_�J��@qJLDXh�� )��:f
��Q�jP�[�|�ux�`���q&�����*&��s��ݔbz|�f�uȷ#�һN)�
���N�y�Τ�@�6�B��s��Ea��fw,y	�qZ9=~+n����`�dc��+Fmݗ�̧��i�^
&�gH������Z���ٱ7��u�ă��ݗ�}t�F)p�� qޏ�i#�IP�;[E{��֣�#���l�Ss�ܚbtN����HtQ�ٚ�sV�cfc�{�@b���q�37���35W��Ed�gw�7@�Xl�P�^1Pc݂�К�v��t�G3+ my�N�p{B��(��������aw�_�Ņ�k�F~���p�w����kŝ�خr~s�џT�|�?�[r�]��g�k����p*��Gmj�3o�ft6�S�Mye���Jm�4����)F�U�t?�D�ҫ�`1ˢ���,���Y�%ؒ'��
��D���gNӦ��䇐<��ߐ��%@z�x9�É�W��	X��:E!����X	�K��<���T3b����Iv�6YNY�w��>��xE��^�wldx��U�֬�َ�^���NH��C\r|�ɨ��p�/��8�,���i��ك�N���d-,z3�cdW�x�.u�k	r��vc��uS��o�m�z!��v�m�ơ�a�&P��P畊��ȋ7_��p�E�V��-[�n��b�)g^�ob��}##��8�w+����P����K�[�˓��~տ�j�g�� �n�*v�:i[��9~?E9]r��jg��s��w!ղ7^9�^����8} ��m��<�����I��P�ي�@�>��.a�9�w��񣞓w�;�>����|3�je�I��������X��i|[�;�&a)�y���T��IZ>���3���m̭I���-	��
?��]�#����;D }�h+pH�<����R����zX��]g����L�������"�6<f*���p�x���{jgv�b���C��c|-7�Sd�!hg�ڣz��	�?xJeИ����'����9t��;:��;B�Nl���v͝�D^�>��{����
��oƩq���!���_�PXPX`Ϊ_=�9.	7�J<�,OFM����K�X���	]����:W�\o5�>s�5mƔjd���a����e��ә扉g@pK�Jn(� �,�T ��T��k$�(���ƺ+�G6(�i��/m�JO�FcR��PO2�&m� ��^�iL�yߖZ��xYqN3z��OK��?��_/<m� `h��+;�X�������6��ta��v�n����O�<W/ۧx�4�B4�C��L�W@��~Of��c�j�eY�M�!D�~���L�\i��x�{ ��е=I��De�B��M,��@!��,�K/r^�e�Uc�,s<%�,C1�*|�8�Q�ˡ�/�����7��m���]i�oΗ�WeiEv�������3ރ��o]�b��|��-
�5��Y�v�p2_~5$��f�`D*��v��
ĮhNav���5�q��W��|xp��<���ɶnam�?�2�k�S~S�1��~H�Nh��<8� �xKzb5�#@`��.e�c׽��3�Y��@��q�U������j}u�_NT���t����6v�̋�Tֽ�H� ��;���i���C��R���7������*{1�gR?�T���w	|3:.�H�pn!5Cm���}�U�`���"*���I60eh���x�d�-p_�k�Qkk���L��,z�À�|�)+׸��8陦�'L���r������2�����F4?��J�$}ƣdr)�V� Y�P6����VIY���+=�/������R/�����
�N�OhޫQ��Y��b����4}�G»g�_����Nc�&�f�c6�u���{3+�e�;D��^�ni�[����N���&�i�n�;�R�����i�3�o��(�g߲jU�-U��)�&����+,�a�vՙ50�yJ�:U�V+�S ��F�J��3CN����q�~T�M���5�5t���GN�#��ﵷ�R��zd�,�=�	ob=aV�Ѿ~������Q����Ky��V�9�)�h�-��[���*T����N5TB#Ww1���_sG�S��ڽ%�k�l��)Y^ZؼF?�)������Ӧ�S=`�ͷ���2
���/8K�Y��t���T߇��	9����%r��\gyRa	5-~�g�f뺱؈|6����~��U8���5�
��Yv�3�.�7��o�l�By�碩�x�1cC��*��YZu�]�M�^&4�yЙ�[�ˆ��⼙�W��!{|�~��w�F,�i"ͦ�x���b�C��L����9�]���ÎÃ=�̲�*�&n��l�RC b��;Ϧ���<�����z	sH����<���e.Wy.E��`�ݼC�3��rQ8�|��p(�سy�W��UY�5E��g�^��ޛ	��^au���C�1��҇��ҧ�Fk��ȧ�{U���3�
(�Ej�X5��o���-�F�VMtz��H��v֫�F�3�02�Zܗ�O�����l��Q,DV��~q��;��Q�+���޵��>�,r���Y��E�Q����+�|5G���YahHFe��ؽ�yO@ᯔ�N���~�5ǏE��b�֩������[jn`-+����i��̴�oz���c�Ԟ/"mf^���P�"CYr)���p��Z8@��Y_�j}����1ۖ��3~H{�p%�u�'߸"%٭ ����Fg*�s+ ����o���4Po5*�-�{���%�;T�C��:�Վ\X�Z/+r�ZO[v;$t}wԾ��B�zf�с*y&=ed����[,Q�+�~U�ٛ0�yC�����	�\�e�_8�&�4a[�C��i���e�z5�7�x�x�E^i���ʋ�����z��n˄g�AU-�7>��~�ִ����~�w���#M���_�_����=U��R���c�˗/p���.Z����h���.�`~�!瑤�+��L�3ʮC2�p�������9O��7������wj�_�Q���`�Ʀ���Z�桏���=C��ژ�{��&ײ M��s��!��l��i2���/PƘvk`�m��qde6�� U��8כϭ{�*�8Qь�%��{��AU�]8L����� ���i�pv_)˚�B�L�bo�N���A1�u�����c�A<�.S��j�W~� ���ݏf�rR�\�t�AV�_�Z�5��v���2��̣���+���-��pƒ��0)�4�������v���Ȫ�>m5�����ؔ�ndb�$x*;�F����b#�u�6�����y9�}Ӱ�u��#5��z��5���/!��G��F�	�(�y��[0͚+�2$|�Ճ��07�~dα�њi�v�3cz�(�1lTU���~\��hE���]��d{j#j\��2Z��#n�����7��%�Ǚ�1,��;�|��ܽ"�s	ѱ/yl�ڣ$�δ;k`�ީ'�}�L5/(�o�׭��|�m4������exA 3���x��c)�~��M��'�J�Ӯ��~lѮ��pF.�ͣ���5��������g)�ɖuF�FL�%��������ઑ���­�{ }�#����.u�lp�GgT�5���ͷW3���a7�P<ϮֹXsh��!<��l�
<�Ӟ�HL$j�m��˹_�_k�N���R,'V;�Z�>^rYW���H{%9��;��|3?js�/P��Iî��[W(�(�S���J7��y�y.m����?آ�3Tu��l�Э��1C�yO5}I~�Ɨb|���0���kS�%�yE�_H!PY�4�K��<��}�X�F�-g���>>���d�o&%��u:�c���00ܚN7���(��ne�{!4mi(B����Q�x���˫����!�اn����j�p,�׈F��2=�سD\ͧ\��	ȣ}��f�ef�&<�{�+��˚cQ�Gs���; y�BV�xz/a�ao����1!�*���i��]��C��Q;,�¾-��/�"�fR~ϰO�qKq8:pppHm�_.�	,�I���~*��
�w^��4^���	Qާ+xZUs�ph��&�g4���ƭҸh�վ�6wUq�BK��b�N�c��4�hb{7a��}�$�"8���9ڝ��!�M����Q��G�MWa��H�}Ij׹杋�����1b�8Z�����v&ȍ4lH�U-���=���?z�W�rO��M|]X�%3��Ny��Wݵ&4����(�WK��w9�N�Y��6Z��66h{|�_�7��p�*�V�?pH�eu�Q���
��:t�Nmo�E�wC�RY�2��x�A�z7��$�L�ݦڣ��
˞���i�i])]�o(�/^��$�o/��@�P/g����K�j�̏'���`����u��[��P��r�r3�a�GO��������U,�z����s�7�_�[���#���}�nC�z"���K�����"��)2�ruq9�a�4��
gŹƽq$�I-W��{�y�kt�<���s����	��υC1�o�!]�n{�x�ϿHxB�~B�!s����u�"��e�WE���5 K�ƽ2=r$�#3[�z�b���[�/÷�W$�w�_�?�D�� cH?c�̈́�|Ľ7�f8���G8!���*}�U˴������ �F��#��5�KT� ��0�[�M�{�b���v%c%1?[G����W#;��Y.����D��WV����8�ǌ�g&I>�F�����|�#
=�}��>�Px�6�r���I��UW�ŵ��m�`S@,/�`�a�sFÛL$!=���j�d-�6-��,{�N�Z~��朑8�	�>��އn^���
ЈX�tAzɐD�;�ӥ5��j���i^�����U��X=;�A�tŲ�0|�����ɕ�tҩ鱎&��#D�*3������r�m!�ӌhmR�2�r���Q�n���&�z�8���sYC���W��4�?˧Zn`/��FE����#|��ǲ*�� zS��	��UIT�Rd��qy���g)DN�l�|),������s2�8���~�X-���ۨ�2BR-�*X5�' ��~IQ4E��e@[�vۻx�F�p��i݄�b-��Ŵ#Q#0�XFuB��7x�F�ū(4���йnl���W�qj�[J�K���`)����HVmR���Bi��wYg��u|7�I�b���j���	s�嬨�Feӟt�e���=�+�0]��2�������1��+Ɲ�8�Ɂԍ
��&���=�̴��ܙ]��&����eJ{�\*���.��
�u��J 9�����O�Ic���#�,����2X�.H�h#R�TJ@��?9N�=@�@�|?�~�2'�?tN�wL:�?��L���/����?��r͉���$Ю[6$���y1�%��;*#�%y8�OtvvRf�/�{�G;I�	�Lʼ�p����кM�^H�<_��4�����y@nͤS
;�0kry/|��T�R�ZT�)R��g粀�XP4�,�/�Q�y�4R���Oؕ��GHX�k�(���ьE��^�����^��}���>���tIΎi+�Jt���**����yc�vH��Pa7A)����.�4zؼ������Ub%����k�45b�$f���hƨ���	�&�����6'zo���ºoؽ�X��zw���V�ʂD��@ᡧkA:=���V�T�m�r��Q[�"����3-QJ`9�~md��(��-�N܇�Wy]�
��q�8�g9�X��K��J���Sؠ��q�F6���Е�Ĥ�ʩ�Ys9��(��c��f��p�����S����x���G.4¬�ʝ���7
a[8�������(]ąi��FS/��}4&�%���7غ���y������}����>�� �93{��{l~B��B���KC���[�w��J��?Nv��]���e���#7���;;f5�N���8u.��ے}��Z��6;���e?�q���*y�@�����,�ٹ?�O:�
�4�����U��tҶ�w�O��1:�խF�2v��2Ig=��5�3����3�ڷ>ӑ�N����}5?�p>L�A��`zҦs�E?��Y����*�Y�9<֭�Y	�{��DU�(ܵ��ƥ��O,�,�9e5,�ݣ*�-�zjLs뇰%{�1��8��@�\G0��D ����,�c��H����љ���#���OoU=�f`���x5�J����>)�`XdL�h��pQʱ	#9� ���y����G�/IX�0-�0�4b�iҶ�y�:NjE�#@�n���Pj>��:8�����C�R_7F1G:�'���q��c�]އc0f�ol��rO������g"�@�V�~ѯ�@�N�����5�t!����A츶�x�_�X^#�vg���N��Sx����ĵKA�J��V;�/��<.�C��n�jfSDa��q��ˌ	��n�}q=����r^(@�O�6O���S߼�w�X=�ܻ��쎗��������������),�q��|�����|�귇�76�Zc<|���T6�� N�D
�Ӆ=.�ݽb�k���^J���N��wL�]�8�El�ͤ7� /��	��"IlzD��;�*���V{'5I��<R��mKY펜�11�\�5؅:�U��g�A�M[%U�x�b�Ҡ% 1D�*x��i�kl���� ;����zN*˳߱�"'؞�$t	�"�9��H�"X4�<�;lD))�b
�v��H�R$�@�E��z���8V22���G�_��*~d�����&��=�#�>�\�z� nn6y�s���N&4��lR�Xٶ���f�`��L#S������͝�:�	���b^��VLk�f�ߌ�.�K�8� [a�=)teh�Y<^{��c,t':�d�K??�,����3�+ߎ���P�C�S,�	P%X�1M�u��
�JJ�ݵ`�������
�ܜ��ސ�BG��d�Ԛ�h\��
�J�(AJ�.����P��J-����cdM+3%�Oxz7�#��.A@�C) `}��S����KG2��І�O�׉\{���ü��X�Ze����c/cl&9�6�]̓Q�x�֎�'?����tҡ"�<"�G
���X{�uϿ ��Y+o�ј���ˈ4���v	�i�n�G*�T߇��]�7��S(�m�\vV6�z�v�D���z�%t� L�@Ø$G8^Ӭܠ�Dk##�>�^�%��PB�oi��ᗯ�,g� ���Dt��i��䘺 }��V��C�P&���:�J���[* �����<��c�</
�.�����s�<��W��Z��@Ŝ�Z�m[捝���Q:�Q����rP{�I6���M��3Rt6I����@�C��]b_��'�n�����;����(s0���2��}��A@d�T���0!�a����/���m���k���P
��&!x��j�/y�{X	 U�<�&�忑�H��ŵ���!��F������1�3�X�x4�qfM_GK4O%����"q�b֬�{ ܙπ������X;����E$���.|�ޢ,��Q�&�?�����-�,�W�
m��f�J��%�������A� �ʸ�����Ԏ�5��;����1G�+���O��6@w�^��+n�Sx������$||WUi�-�2��B����������[?���)XXx����R( ֿ#&FNA瘉�=Ӕ����s����b��V~8��R,p.��%h�����wP(͛�(��#����C�W�W���R:#FN��w�(���c�Ai�n[ʭ�`i����8Mτ�H옒�ŕ "��p'OFY9�]� �&� ��C\�81|h�/n��h�L`�Tq�ډ��Q�6*Q���X�N�˼���{��!���$�
o 4bDqX��b6���&t����j�����@�����œӜ�p�2ϬL��[��R�5$�~�nq�*e��8JӐ24.ƫ��.�=�����6gicT��7�&R���#b�y���q�W�_wPsQ�«w�J�E�X�>'�k��h^�¨�_��)?�D!��ҍQzS=z!�a�agqm�3T��F2������Cb&Q��(?���xh#[Ii�������i(�Q{~�����P����"Aa�1fI z�~���X�w�#	{�@h��2���@��lҹ��ߔ&><��蟾��'r������������R�ܠZ�x)�Ƥ�Y㽔��_�G�Y�"���^�1���DJ��Hq:zȻ�� &�.
*ם��i1OzQE"E���A�IpY�c}��X�Z���~��?&EJ�>����@)�,ZG��uH���/r�l�p ��&�n�^�KHK�;���r��ֆ^e0������J�1�g�ֈ��:�.��s(@�>�_ݓ�֎�j�MYY�HA�h���8�@�95��C$����&z6zsg�9xD^���V�)3�B8��6�i�6��O֠,�
�I�3�u|��E{�B[�W��0HY�ؒ�4s��a�?�B�2��5C��~�︘����F'2c�4�Q� LL��f�O�|��К��ߕ���S�q����A�֖J*s_�����ή���/��q�|
!�8!���7��Fl�N���h��d��9�i"F�8��l"�O|�@��ǉ))�4���cr�'݆9E��\\��Rs�w�%�X&.8�AF�7��l�@�+H��$V`I��}F]�S�*a�������l.u�vGLEh�)g��4h��Il����*V�����嶸��mY�\��q`74��J����b䨐�BZ���{�۝d�H����xZԉ�)����^�Y�h�S�3�%6�$s�4Vp��cF԰����3C�����C�
�Q)�]�̃�&�$ְ��P�@�l+��=�tLS̲X#9�2�������Ñ����eܚw���ʣ#C�}]8xaIgLqqJ@>;n-���y7*��:�̱yd!PM|mB&]� `���`G�C�N�-c��~>	Ε���h���Ƿv4��6�u� #�0�o8��O�:s�üm��g����w�$I6�>b��+����.��Kj�O&6�j��u�xh��W�D�wD�~�H�K���/�i�i�'W�4w��_�"|N�JD��$^ב&�����cM��']�ƕ5�Q�$�h�X3��Yْ���P~��_	�ڗ�XD�[DQ�A1H���B�.2�Y���8dVjBY)���(��;΄B(#�����eZJ��\�d�uW+��&��:tє쪟�'81>�ȕ�f0}c�a<�A����4�Ԉ����-\eG��	B�Dmr:�?#�txHߧʃ����d�>3̒�}[2rk�׌��O*j7Ӣ����ݬ#o�:�}�#3��H*��+i���X{u	<�^U�u*H�^�"c0��>BS`���u	E�?�G�C�s��bؑ�2�}���V�����h8Ξ��S�ne�x��P�Q�D-!�Rq�jo�����b�p�jͮ�Ei��w�����c�P~
���@��	c�A�t[���OO΍���ќ��I�l��A6�DZ�!�Y���o�W%�^�q�S>�UP�Y�3a=��a~���Ll��F�i�Y��q�@ʲ�S9cd�jE"�{�d�������?Z�l�.L*MD�J�"1��a���ϟ��۟���@]�/S�g!�o�'`��E�����	����YD�R����V�v�`!�_����B�*Sf�[����~_��`x�[
iK_u�3sfC�b�qE�r!֝���("�x�ܕ]��U�X���i��T]}��4�{�����'ͷ�E�KV53���]9j��z��1C���ڧX��Wg�01�@�����3��J`-в`<x����蹘�p��DDz�������3�Ëv�l��D�jwW�f�����)��O����Q��J�h�_���=1�sX/5���M����An:FW@�_�3�0�+����rS�� Mo��ܠi����W-!:�b�+��	����{���2�L������Ţ�8�'���B�k؃o_�H�(<E�2�� ��oA9�m��}�b��*�0�i$\N(�-�O&,�p��{�'����>��"�4��e�y��qK;�k��k;\��YI��hA���c:�ތ����3�I�y��e	^��P68!!ÅE!K�G���lq�0t7&U�q�E\�Z;\s*g�(��{�JH��R*���4*Ϫ���ҫkφj�}�C�W��0Hm\�����t�6������Xk�:�����
��A œL)t��`����$`�8�V;�*6��&I�.\�* RG�=�4-��p���iie��V�@��59���������(zp�DB#K�mڃ�)��r����x�v�,Q��m����#Y��
j?y� ]Z���m��1�x1���}m��e�I�(�Qq	�� `����!x����_>����GE$�4� �*�-Ǧ��8[ �������*��ρ$��M�p(#�b��?94}�T�k��R(��l�ڍ6>�'�=�%�8(���B���/�TH��f�-��	+����]	ә�W�ĸn_����9 ��0ړff@lvT��r��Ǐ��FӇ?I��V�XCU)cPTz�r/f3s�b�wi7 �[g"b<��x��Pn+g�;��<2�ˬ��Ow�t
��d�`�	.j�C�4+��M~;���eM1���.��E2�ӝ�ů�y��~�r��;`R���pr�3yF�w��c�I,ǈ��,�YTB�݀dl���!*�/�<v"����F"cU�����Xz��CM��+��1E��n"���L��Č�-^>�?P�2Nγ�Nn����@���x��>���>��q�|@��̋ߦ 
��l��\��C�8Z���#�=���ȧ,Z����Q���T�]L	WW�2�G��m�VPf��B�y�O��G���Z:��'>,�W�D<Bd�<��6k�4w���/Z	� oΥBd��#���0�iuh��H��'��s.28����0����9�b�E�7��r8R�S�y��Q,`G�?���0��fT��k�W�:�Tϖ�8�Z � �M�
���j9�;��_ߒ]�F��(�х��+�h����¹��1[K��?r��ЇGn7�炽�<E�d$~�zZȀ��c2���M�{�
�򣇪��T��	%?t��Nﵗ���� 6��p`��)�;�+@�u!�%�Z����ҏ����廿�!ߡ�h9�.ڸ'��2ȅ'&�����f�����% �b��s�lC�6��D��?N���^=��k�0-R���o�o���䲙1�-(T�8���QO�Cyw�˰1��>�{�9sH�(ð�^���Qs\-�w��z)Q�'��H�	�Z�:�� a��_�������Y��v��C�'�u�h+4���a_I�z�d�B	kZ
���v�r�jZ��4�&��K�gb n���eऌ$HH�@,�Q�j�ʤ�Bo (��rns5_�9(赁��`�8p�E"�~I6��{zo:�����jydW.W��������Yx�

k����`��TI���r*�%��9B�	�X}�s�PX�2?����
Zj�jpQp���+�����~�A3��!%�7X�U�S_�iMRe<I�Y�L��p�^�
kzm�ߙ'��Я+#)M��D�Y9���Q�Q���ʩ�y�s��߸aP_�g�؈K�-��Ӛ�XЈ��M����G�l6޶��`^G�I��z��}��1㙨�|&�j(�?�w<���o���qdܙG���gf���df��C��9{e�^��d&�EQ�B!EB��������>_����~mtW�fo��.z��k����̯B���|P��š䒕j<OV�u�cJ��5lZ�羬�M&��̈́_jk҈�x]=ͬU��7���mepQ(�~ƫ�/�)ZZ�|Zv*�-�y���$|�/�'�%1�b��07�~�4�S��UiV�
�G��w�i)���ç �d��~�z��u�(��Cr�I��J�?����(��ܔ�jr�}ж�˃�x_���AYU���,:�����Uq�h9�}���pG��i��5�g_F5���2fu-#�k��^����蠜�S���`:�zpMnQZܽm���/�!�<jt����{CP�y���k�x[ƀ��C�ƒm�߄;,@Z�]Fҗ�,�'���w�ݠ�JN��fu�m[����_�Y�u���ί�UpW�����9N�e�?p��$E�6��A���Yqد�kXqC?k%^�7&ގ#P�1�G���q�xn���e���iᆿ�@Bzr���L��\'g'��cؑ��w�+��l�9�� @�R��[��D̑��d��Z�ƿ��vLj��q�q(����$J��nw�9�z�us�c�jR$�M8x�.�^�?��ti�y<S==
�5���Ȳ+�6󉊽�S?Tג��RH����3ahC��,��:���(M�@�.��ý�\w��,���=r\�.=�����6Ki@�*ۻߴ���Dz������Ksf���݋h����0�ۼ>�+�� V�?k�y�(3���o`��5�#�v@����mY
�G��)��1y���0��<���$ �RxD�oC��M*X*htJ(�R�:�~���db�p�4;C!�M�l�V��ȵI����܍��〘̆<�{m헉��ÇE�QClO�;怓V�A�{�ٻ7��	�����yaW
EPB�I������_��a��FsM ���~G|�8���{T�K�c 3Lb[�
�����<of}vI�xզ]��Qs�rb^��n#�]g����HL�L�����roj�y�}{�q��q�Z[�u��� Ԯ�@â�񭩢�����fp���~�G�-)/���{-X����O!�{�����qf�!��5�Ϲ���b����?�mB�j}C��EV,>;�~v;	��@��B-A�U�kM�;��z�	@l����kM]߿帆<.�2_��z4$�'���Z��*��[��?|���n?��*�
Id�'��5��*��iҾFW��&�:	/�NV�N��`�i�2�Ľ{��ʉy�FS����V���%O����8 ?�̕�Z�������Y�/���h�m�`�R�t�9�´ޥܮ�a�)��K�GE����� ���@��㎿����b�a-LA�I|DK�����7����̓�� OAC���$3z�t���y�$�?4+�UY���zʼ��3���ၪ@l>(�<�V�Q�/)ˋ�3Mk� �z��� �()`v���R�O�ӗ��m�)O�,S����>j�'��s���>?V\q�.�X��v�R����t�շ��_�R�i��Ŕ�3К!�rʑ�).��5���S�_�2n8�Y�]���X�bT��":b<���O4 \2��ţo��� �����cg���U?
��)l�Asm�Rw�Z�L�w�s��i��2�����FK���Mʿ�xE�L��V�=m��/E�a�%�nݯaA�ap������E)��2�W�Χҵ���:�E�s�)����>���D�m�L!T!�.j�a�æ��e�S37�XC�.��k�˚F9��ë�J<�hgŕ(���$��e�y���
<D�u�ҭ&��hQ%�
6�_%�u6�[6V�2�G4���V���L������Z?�SL8g!�qA}	cuO����-2�BΒ,��d�{WoD����/�^@�%o5x���:���4eX�M*�1�㩨x�b��H�)IN�Q�ƚybS�?!I%@��Fq��>:�-������k�S\��];�0K�Ѡ�CN�3�*"�6O��C��+%�TI���/��kf�_c;NY�+h�|jv�l�j��o�UV�ߺ���˞ٲ*�߼=|�#!n~�-�8����Qג���7`��J�2��u�JD��*%��72���cl��#��w����e�����"�}�d�|�U!&J$�d�-�N-&)��Y����$;Γr��>��f�vgĩv�,��f��2����Լ�pq�j���?�=����.}�ڋv�K�Z��ߕ5MO�~���r�o���C`y%����S���ͨe=nn M_>z�(7��Y,�N�����C���4kZ2C-�G�#�S�����ox.�����H�I������EA��&�9�d�Y��uE[OK	-�{q}.����5�p���H3?�`�wѾ�H��'~�bld�&=�|�߶���=`a�N7iǉb�'��`��;`SI�|��P������NK�zχX��&�o�	�x��o��M�۞��h^�fv��j�'�f �����G�҈Y�{%&�uZ�/��}]]F��c��uϐE���)�j�P���"J�S�o�������8ޝ05�����泥t#����D��WÄn��o��/\�@>��\r��eT��?�>F?h�q�^nna(4-)�֣	3fM��O�KS�sq?a���Tf��V_j,6N����}��-���a�`ƍ�6���e\� S�cM�ک��QP�}���G�l����&�����D�A������we�.Զ)�10p&�O 1��W9�c^���};�ɏ�4���k��F�@����`���X��-��؍X��p)��������7"�Q�iU��	�\�b�;ɭ�A��e���������)N�gT�3>�4��M�Y�p�U�J���N-�*��m���=�ۼ�{7A�0�6h�p�q'q�[�0GL�?��b���-��X�9!�Β�e�oϦ��B�ݍ��U��.��%�ꢅ�f1_�+E��c�z�쟓f���-�b��yհ�A+��3�9рcV�5�]�����������������g�#�xq�bt�HI� ����{M�� �1�N:
%��[�%�2���q�7��)@8�����i)��򸢆�C�I!���	��Ȏ_fM/�����D0���@���S^O��T�h!�٪�H�#�7�0y=��9��wsՖ�����B��hr�s��C��>a�%԰���R�B�3��|�����v�N7-j��(��[EO�!]EBQ����וv�Ԍ��|�ʺ-�9�Zה�z�T�	k����L��^�Z�8�������Ǎ,�k�i~��Z5"`�<��+@g� �ޖދ���I�(3Λ5_)�W��A�x�G�c�i�=}ޖ���u3��L�M�I�$�%{.�;/n�qv�́
3a_��4���S���g=.��t�z�#�B��$�b�T\Q��Ld��@zj����ۼT�� ��!+�f\2���剦�'@aw%޳͒�x%p�!��^��M��DDde�,}g��j>.�a8�iS)��L�S)5:���p!�w	���H�H�Xg@�<�d�J�oj�\�q�#��)!�$�y�	��sjf����	���>��8o�u�;'C1-+
uԗi��$�ޟ�L�Ѭ�v^B��g�h!�jMqV�kN�eZr.��"�'^v�@�Wq���Ü��2��p��
q��@|�D�T��퇥�j19u-�򴻎��Z����/�?-��"�f	��NΛ^��<J�:y���A<aC$���V�v/����{���ŐB�LX޿E���~�����pf��$.�fYv�����n��>ӯ+�(b�@4<�IR"�!��S��d�H�±� .��y��f��|/u�Ҕ��^�{A�6��xZ��*�����Ҳ�P;Kv�h ��9u�"����׳
}Y�7�-a�$hfu�>��B)I�*�<�H�Q?�O���B�Q�Y}ژ�\I�l�P_�Tqd�5�6�N��I����G�'�zۡ6��Z��c��_m�;1�U��}�ͼ{��]�F�ƪb��߳'֯�ķ��?��	����ԙ���&~Ǭ+i�����܎��C��ig�N�l���_�.�Ϡ*}�ׄ�Z���d�
;��������t�?v[<D̗M�j-��(�;�J)��(	����%Q*�}�'�F~�z��($h���o���p�
=�a�
i7��V԰:E;�n�,,���>	��a9d���q�D�dF*����
��쫣��1ǂ�Vք[5��'<-�0����y��OB;�.�{��'vY\C��>�'��xgP�K�"�>��߀u<�Xd����6�A�X\9_Hڬ��v������ix��Y�,�G5�7��l�kj_���c�u��s7�vG�7q��g�<*M�������a����0��i�.v�Ɣ�|瓕�e��Ѩ����ť�!��a˳�,�If �z�e?� v�O&"���ɅT��,w ���ހm8��/�w�4���G;ǯ6�	�_�i0����]�q~S�C��5+�2��qIj��7AU�~��~���OO��5�8P����;7������<�f3�yL��Z�,�m��m)�A�Q��u�lWP$@�S���\�g)�v2�<�f�F�T��l�ԜtdxsP�7��0v�Y�v��ͦ�pf�������Q��_�鋛;�����|��La���r57WU�C��&���w{L��@���o}t�:�Z��QL�|R�y��o�K;њ�cZ~c;�:ED�q\@_�+������s��q3�Tl�W��   ��$�%��c���[��'��������<�"'�q������c��ݴxM (>���B-�|��E�X�^�`VÍ][�e_s�]��^v��q��0�l!���~l��tu��*G�D>1c[S,s���M"�m�����z��f�;B(�-j��6�6��j�0 �[)��-5����B�&[��OWck�^�����s���D��n���;�Y�5#={$~�ڻ%�,9��O3���󳨜l�����	Wr��o�U^�lͰ�J�������V��a�eh��ǵ�ϼ\��ʼ,o.�=L5�W�W�A�aC��i=?��*�{8{v�#�q��? :*O��f��kY���b勂���`��[`�DC��J�t\ݰ�xTq�^�z���K��`��~�W��I�NzK2�h�J)�Ѽ0*D̂�&+������'���~��m��4w#��d`�JfTX^bX-��K���P��e���7��
߰��NJ�ç��IҘ5Hp���qn�rAni7؝x�կ�RM;4q�L��)e�SQ�=T��}e���F��kj6�Ӭ?�v��曚-j>��o�������"��o�W0�G�7Є`'��'"�||��(���H$�� ��D�?��-R�`�eC���rY��t�L�A�[���4"�3ر�q!��U�fm?�A��i�M�k��R-�&��4M��GV���R(Y�B���":�g���bj�,^7I��͆��>z�}h�)\�(�m�JV�BC+��D{��$.������?�n�b�mm
ŀ��T jY�\��N�0h��o?�]��d䰩*��9���oXlӒY��uf��g��~����mx}�Ag����χ��w�v�f�Iz	��bD&����n�
Ґl�v�<���Q��%���9�z&CE@��XhK)N�޾�(`�y}3�Uw��D�3������v,gQ]�=��������K��9[�]kl0��o@z��~�~���������*��/.���0T�%դB�=���a����~���<v�|R��_z�C�c��,�v9�1�%��1�y;�W3�I��UW�+�G�ͩVG��둙�:�:-��a�a>�	 ��[��o`�`��HIL��=�eNe��\������l��8_��b��~I���_� �Z��)b�r�:��
=�����K��ZB�Ȓ7�c��,|ɜ8]ŋP��r�1�����&���S�"�yw��hj�daY4��"ru�N'�Iޯ�r�w�H�<5�����L�d2}'��I^��+�kf�H���s�m�.��o�)�;�[1V(�R-<_<y�>lvg��ʼ����-m���$j~5�h�e�i��b�'�;�G\V��J�a�g?6�Y!�B�]�+�)��Ev~����BE�u:{�y{�'$��q��zI�,����y�e��#�Y���> �0LR_����'$?U>�l��ڃY)v��@�Y��m���0����ם8��m����>y~�z�vEB%����	�nx<�O|�A�Y��f��,�}�S�?��٘��"��d�N�'q��v�l� �n8�<��Fs]�
W��o6���aE��KK�}�;J��gY�D��".T��Ӵ�d�-��\B_oS%. C\ķ�� ���8ξ:f�i�x�*	�(B�I�57���sL��p��y�,�:e-�$�f�t�T`���z`�ҍ�wʜ��=͡���h'Fb䄍�F�jьϳҗYI��!.�����*H���c>W�u��S(��a�F���C��֔`�0ñ�����ӑ=a;�6����= e��iB� Tj$nbsڴ������%���@����;��Ag\�  ~sЖ"P���5�	&%��0~Т�z���1�gΓ�X�頢3��0K��#�\�4�8u*h�xo��υ˼+�~EK�ij��|e¤����꠵�t����{��ϙ�@p'̿�o�[b��:R�`�',3(e��<��1��{%ܙ�k��ELR��ß�<��T�O��0]�:D?��}q Ђ��5e�`TҬ��v'�|�
1�L%
�>����U0P>�.�?#�2/-�� dY�8��(�+�{�D��u�y��"�i䄐]Q_H� �,`w����q�&C����}�v�q�-Cn�V/�B���smF�8	�Z�ԴB�V��$c_5J9��bɁO���6�^/����v�F��(�R@[^��N�ߡ����]�i�5�.>�fy��k����&�D�xKP���� �!&59�y^"�kN�r۔[ f3��zQd�r5�0��#qSD�N���T�|WM�hw�W��I*�S1����n�M�D�G�<��s�*�l���;3Y��R?�[�SN�טc�fjsF��K_����XL�-�W���-���������2��0��&ζ�0��/�Ω�q�w*��m㪪�:l���4qc�(�ےOv�R�h�XOE����40�ҏV�
���l\R5�1i�0f�t��)hG)������:D���J܃I=�5*b�2q{*!|ȀdFq3��i��|,����d��y���F˰��S�&ʿk}�<��MaB6%�)��dj�����Po�`�ti�u�*a'Z��-2Qa�t&-东�g�h$W�֐q�e�$>��[��u�������]�͢8��
s��q���X�#n���:3���Ïgv��O�B�y4������i&���q��x�b|W�K1�,��{D�A�����nY��wy�z?��<�l����T���j��p�2y*ش"l�bn��T���|���s,����zP���&>fQX�>l�=o�
�W�ʟc,Ƽ�$6J�M�f�S��L2�ɮ�:�)��.�g���'K�"Qq���N�@��t�Z�3����3#XAE�̩�2���8Ђ��;���a���c�z$�(h.�3�*X�� ���ǵb��ͥj{��YB܄;���=���l��*z��_}��l�Yf��:��y�P
I��rā�5r��W�3e�b�qfn7�����WR戚�t7G�FKu���c��:�7���w�z^M�z��W��m���d���.bf�P�R-���6����� ��{6�^�5��ad� ��"d"���P�Jt�'�	�C�eƴ8�<.�X�-���;%Q�/�3�j��힦O�R 	�WV�X g�y����>��57�.9V�U�ڰ!��m}��<������&s���h���8����T��l,�k�[]����65y���.7N�"���ǌ�l]t�A^��O��n�,�r�>ߢA'\]w����;���fĝ1tAG7�?����WQ.���*L���ߓ�g����_Q�@]u��*	4Z�`G�cج����v7[����UtY�-��LR����'�6����D�h�k��.JI|Ը���
޴}aY��5=  �m��&�_K|#y�l3.)�:�y�JQ0�-�C��><B�{�D�R���j�m5}�0��scZ�#{[I����\��~F����� ����?�L�N-#=n/?��'��C�׸}���O>�^J�^�̏ �DcFi
o�9=K[�nÙy*-ϧ=�چY��V��y�B���⿺Uu�=���m(�/�^���h�h��f�}�	a�ZY�NZJ��IV��J[���Kӣ���N4��rߺ$��~	�$����r��p���in]<����8�֦�)*��\VR'-ui=�0̚|��=3��n�7e�&�F��um�>��9�	aA`f����t��Z��%�jfL@�| ]Dx@V��qN�/GL�:�؟)6թo��|ߺs� ���ڧJM��z�eڢ̗�>h�}�9��-KoyY�r�ڭ��ۡ�ִw�XTΪ-�˲S"���K�T����`:X�(��f���0� (����[��A���nQ ���X������P�af�>��Rvo��u���RE���!�e
P�m�)��#kp����Q(<��S ��wϟ�f!m3w5dy��T�fN.�[��Z���l�*�Zx�$/��mT�C6��+���,zP�>Iÿ@����Eo=�4�a��r5�+���)d�I)�a����|��K��l1�w�'C�?}�$q���a�VZ9FD����5�x��R���;lSZ� 5�M;`�e�o����܎�CL�3p������ =�[J����T�V1��ew�Ǽ�?\fkg vrq�2I�F�����7>6TXe��k�_��yxX���C�s��U�DM(
�7��3��,r�ˡt����~Fcv�0�� DA��Q�b�شN��n�s8��^~g�R-c�~�lsB�7O���>��L
��.����	�G��X�"�"MxUa^R����=1q�(���5�Ώ�|�m��T�j���;ɸ� &������#4��y>h��CNHa{�Td|�d�`u�G_}�8)�ְ�V ���	�� �a���p��"P�;�+�1~u�1���1F$wj8J���ZEH]g�;�R�o�j�Ѡ�/���и=�4cO��8G��#����y~\	+Wh��=��6��!Ζ6�e�0��g����e�h�l!���">u_��BBM���\�
cv��T=��j	��׫
���Й�Z�F��U	�h�f�1��쁿L�nC�h=���Pĉ��7�&U|9e��¡�})��jŎ� U���H�p2sU27[K9��K��
���+�J����:� #?����0c�'�'/���������b:�7KŨ�]M��/����������w��fd[&���v�����yb��V�Q5�hr,:��y�U�c�UskVG:.ZkV����?�|�q��9��e���V�En��M��3}uF>�_%��wo��~ \E��������L��J  F�T����^6bP���VX��1��B��1_Uó��.>�(W5�W���"t�e����S��'�#_���l^��tO��Z�9�ь��.��'�bV_�sw�����(��]�T��^���{�9����xC7`j[�J�o^ͽ:'��}���#2Q���"E���Oy��N]�5�r���1w��u�����9��훛��K�
7��F�<��o����������$������E��o^\��#�^hy���Z,]7�y�ߑè��z}~/(��|pa��uB�5��*ޜ�
G�yG�&A ��^�����F�m�q@�ݤ��	�U���'���<FU�3�$+�.��@#A��Fe'��8@�ݠV���:W�2���c&<<� ��Jŕ�c,��#{��p/�h��`�0�aB����ǃ�+t����^����F�W��p/�T��s+Qwq)$��_�@�`(���>����Ŗ����R@�#����9���u��~���Ã���:��ˏ��n�{g�U$(ޡg��[D^V^��fY�4��I�:��h�+���t��5\:+L<�M��7�x��r�� *2��Ue��7��t�y��{��^ư�^���6�Ek6�[NO4j��9!&/����s�A.n���ɸ$5P/P��Ƴ�X��N��g"�@kv���b����d�o�V�#n���9Z=#0\�>n�N3��>Ҋ�,�{xd=�d�`��ݤ^��D��*,'kZB1%���l(�F���`��g�N��
̜B�d*��ZUb)K�m�9������f3�$��X��Gw�W"�e��V���7�>�S���>���9Nޜp�(`f_&�:'T8�,z��sx(�}yB�������y��� �Q� Νg*��*�v��uZR[�
l�n��O��� 5f�&8AI6{U0/�IG��n���zPV�,t�LI�%�2z�˪Iv�84i�[�uɢ�u'f���kB��UQ��>d�IL����kь��i�w�1�;��#�(��ötS	�Kbv�%<㝺�`.ƪ�7N�uv<@�|�f��p9��M{N����y� ՟�}:|����;z�'�K�`�W�Kf�4�h��ȫ����B>�ݖM����.�e_o��#�}ԂC�ReC�ޤw2K�T/�Ct��LK��`�+ q��cE�C����zg_7T�̣W�t��t�I+Y�(��#�8�j��yPg��۾�<�mC�r��p�W]�'�'�M��W�C�J��dn�j�;��Pš��������b�f�E���8���z�ZֱCq/��/Y`Zؕ��b����w��[�h��s����h@p#�5������W4>p�~��"��;l�U$�K�2�r�mҍc�3VYr���mJ�2gˇ�	G�Y��`إ|Z�T��Dg`�,HA��z�+�6����;�&^�܍5KL����]<Pag�k@I&���B?.�ae%�������K
���t�yyh�׃��{���SiAQ�\������/[��.~w�e�D��/Da�:���U�[���H��lإR�6ab���$���ǰhwRб�t���y+A�9(7I�}Q/H��n.�׸��Z��-�S^0�W�v���u�z�8�����o�--�rڭ}�	�3��00Yr������|��8D�-m�g<���r��e��Ƭ"SVKB��S]�7�]���b��ܫ�1�˼�i����{��+�R@�������|�n���D��L���=���D�-V��I�2�F+�J�iN̓G��Lo]`0je��W3KX�^���ac���3H�?\,�j^�n%��q?�ߪu2u�%���t��9q��U^շ�
,�\���2�I�p�;�.��m�(�ZV~�wj帯-��5�0uUu�a�_z'�K�"����rE L�ykL�V�w�v�09eE����LF�P�]���� �b�T�IZi�q�ϟLhqT�-���\VP�x�ۯ�O=be(T����x�K)��&�F��mZs
'\)����</�ĉUz?,=b�Oj��}��s79�UaDJ#S�(n�ӣ<7K�U���ԙ'}G�C��Z�|T�7���|�b��`>	R���Nk�+F\zD��4���?D3���i��zĽiʛ��gz&yQ"�| s�*������W<@����I��".}�!����]?�_Y�i ��C�C5�:�}%�Ȟ�\��u?i�[zq��]�V�����C���,���t+�:���RNf�m��(>�8���<b�\�=� K�͝l�
o���| �!{�LG|�0;sd�vD�BJo&<R+32Cp�ک᜙i�a� Hq��<ŕ���䆢OQ�V�|SJ $�r�b��`K5D�\�)����:��
���W��[}t`�W|�_�����_�J���HѰ���Z�ө���UQ�D�1��c��'���F�e-Z[�j|��Ώ�3�
d��ŷ�_��|z�E�U���b��8Х)�|KO�*�Tg��*_�bʡ�ʙ�YK�V;�X�ڏE��8 �������ڪ�/���&jC����U?����3?:��t(&��'��\��%A�����q�K�-��M�4�(�*����Ŝ_
_��cf�j�2�#�r\��z�ě?�"%�ʰr���{|�e�U:2[w�s��K*������q]���,���\1�/w�l����<��D9�qqE��5�?h��L�����W���/1s�5�����eA@��H�5 ���S̘�n��0N;cZ�|���o���-�,x��N{��B��us���4���x$J@�p[&:��B���3��M<!a_�=����$U|P�pr�s���d���6��h�?���e�['\���d���j-/���끜�$�{�Ct�9t�Ȕ.	�v����w���.��(x�T���F��=b�z���E��l�mW����gRM؁+���1'B����Mv�����BH����z�����rq,f�#x�ؽR	��X��Z/���hBn����|"� 
��y���Ina�ڰ6����A�ʘ�}��(�~�(?���W�zb�"���g����~���UsN���b~	I�3G�l�˚�����0���|CL�"=���)-�BM.�o���7vP�2	���JB%Ԃ8�݂�J��T�¥[򼈽ε�2Ï�Xjn�~iz���ۋ�����|~K1q��^��H<��c~���T=	�!�9z�i��D�?��͏1�<��w��+J
m��#r����
6�������
ya&��QF�uK�)��Q<C�`�t���B�@80ߣ�-~,Ĕ��ԗo��E�������n��C�&[���'�i���RC��L{9�'cd�A�L�7YL��Z�3~\Ql�Y���Y/�#�OV��M��G$�L�]ٹS������yU����d�P�|�&�T�ʲm��N�ˏ�V�<>��+�O׬U�9�jIM���%���������C#����eۇ=�v���Rj��.o�XIa��>�@7��t�H���M����������rT�TB��<�x��W3�@�@�|~�٬iE�����G��O8��,^��J>h<��i�E��U��U Ŭo�i΅�C�٪��؆�R��� �F[D񊍄$_�jf��8�шZXB����S�1��Y��+�Y���	M�L��,'���J���c�R�n��j�jҶ@	���^�/�Ʋ,8_cPgP�J���0U�D�s+�Z ��s����s�)����{�5�$;"m�-�|σ���X�,�(��^x<Ѵ�dzbտ�����������t�BRiJ�$Y�~�y���:C�h��8!��&-�^)7@�t׍�a��U�W1�`���B���hT>�f-�Bi�j��`V,�y%�3�E����X	�  �27x>3���*�D��
%F�K����@Ȅ~�$�.`���Q��_l��r-����<�o��h.�zQ"@���U�Ʉ��*���g�y��+J���$�N�^�]l��I�I1e�R{m$���M�B�T(���A�ڌ�I��%}�-�7��{>&��6��5��鬴�7����cN�Q��#��Ե�]}�ԏ�+���"ۆ��L4�3�<�ذ1�R��8�>��I��K*T��U,d��N��L2~Pj$|���[�p#p�O��rA��_;���.WIc�1TRa���L%�!���-#��V8F��+�I�ɫH�]�v�@eA��`e�3e:�Ԫݞ�Hh�Ľf4X�08R�󦝭|� ^Q� {-��}��m�ڍ��oL�ۅ�T�`���k�N�/R>R���.Ǻ�����8���
�-L>J�|�_sPf�������������$l���kpL����G�>+?+���3f������N��1jY�x.�wEx�b�B�ʌ�v�&}�zjAf>����%��JW����,"�O�'5�$�Q�t���m�Go�u�%_G�1��5	p���]_�r1f�|�k��F�����i��Z\���z����+by͉W��o��G�&�_�+ш�W�dx)�u��V�kK]Y�h���-�1��c��G~�����R5ko.|9q3W%�^yw���6��֊�])��*����6�l���X��`�sh+�����l'.w�>��I���!˱*���o��zy_��=��f
&���|���cn3���zI���[Wq_~�L�<��Y�һ�o��>j]ƶX
�x#��Ɍ�PmO�C}�w�mg�̷�ǃ������8}o�^��1�����)���"���3�G��Ul�jfS�m�:sj=z������<!�����L�'�y���Ԋu�{����[�L��s��	߄���n����i�TP�s�<å���M��y�8�_�����������И�7��eA����3UE,�GWgu49��]s��z��GV=nh��Qe���;����M��}�;�5-���5#:(>�����qW�G?V���s�h8�껮�� M��"�:N�
���<Y������� pm^�
q��s�����7l��.�~؅��r��aK�z������z�O����<~�?z�U�u@p�|���l�A��7+�wg$n�<	��N�^�K6�-�,���@�Mh���W� �J8/��h����y�W5G��,g6��ש�įA:F8Ϟ�\��p�C�M���x�C̅ճ���f��t�f��}8@Z���Dsq\O��µ����(�����[-v��e��\�@>�@Y�p|�� �������4 �?�ﶭ� ޒ��pe�g�w���[�@���d��)�_���IF�C�A9��+q{99�%S���M#����e;a,|l�8��%�=Њ_㏻�w_l�M6Y�hx6���1㹺���1)�cS�Ap`i0��u*_9x��������
��������p��w���/C^�G=��`:�� ���|-��6ؚ���0Uɳ�Ӿ����w���`=��Ȼ�\�� 1��E�d1��<4巧 6��������'�t�X5�#��� @7 �c3�߶}���tK/%Y�n���z�j��"��0�v���;0HOըq��2	��D��Ӹ����)@�Ӈ�I�����e��Y��=�8�[Y���'�yh�{�m  ���ZjRz�_��c����<�> 6�j%�Pc�]��_��g ��FN���~���[ݪc�Ԉ���}�4$67o3�~z
�@}��� �:���z������n#ߪe�� ٛ�{Y�9g�v%��J#���x#�㖐�`��sw��c���N�1:��O�N���qO�X*�³��X&07d���>D� H
�RY�� ��83���Y}o8����:� ���+g读v�K
d�\{ ��ⷺ\xK
�31��qKF�.t���lN$�e<I`ġGI!z�l���D��5$��GT�y[3�l�z�" ���<�y��q <c��g �8�HI�6G�}o��̯�e��rtZ�^6,@D>��<�Kߚ��N��.F++�{lfg��}��b��5F����^���J�6�&�V��?c�|�(V�<��>�#8�M���ۼRbh�����md^���?�]��\����3Y咔5����
+]������F6α��ː��4\3����zP�U�i8��CB�to�P�Ö���B��^?C���[��4��r��5d��k�9D�<��X`�z|駹��!��]~�i��Fh~qvQ	��8� �� >��L���4NJ�`$��d�@Ř�}�5iE=�-�%vY7a�C�R4S��ލ� ��/c��Qu�o�MVP��,�qax������q�AM0ѻOB���B7@I�%4��B/� RB�
�H	��	-)�JSA�ޛ���(E��g�{wv���~�3{�9ϗ��}���lꂌr���g#P��ϛk1>�396g*u�-��f����B�WnK�^	O�8�}r�J+�2;��s��F3�ѐ��_������q濪�+��I��_��"���+�~z�ɀ=1�a�Zd������x�bq�A�Of˙���T�Z�2�VA�33����S��";� ��'�P��S�j�w��E)�~���Y�զ�h�}K���Ql�����KTp î,��j���LS-��#2>މ����Z%��-��p��`h���f�Ȩm`�&����ՀTG]�~�s��N2B`�D��]��r�Dj�ߞ.*�9@������K��<}��k�9r|?���]6!/���B�|�̾?�?��@�iuJ�Ɂ�ElP�tj�!Ⱥ��u\O�`��w��P�`��5w��|r���تi��Pȏ-������,ػ�ʰ%G9�~��z��O�)���W@����l�Ox�w��Z���p�Ԍ"`g@HE�;�5�Q���4L���@R�j_|�};����.�d� ��1$?޹�b2����Zŉ�CsCf��2�KF=�x����UIE�0�p	�p�i9�����qh@BK���-�H���Y`�J#�7����r@_ t=	`�-�左dJN��$ǁ��K[�{B��,������q�Q�,�5_SK����&e!L���T홄X�������lp��}�8>D6�ط��,��WL���4��彩Z�d����~E������.(���̤�C�E��[�_��	���3`J-�����V�-���J2�H@�i�tǉ�@<E|�!�.��C}�q>�:�R>y�}P�U-�܀�H P���r�����'n �|�,qi�U�+�x����
�SUP;쿩Q�F��H�?�_m���iI�L�5+r�
Pr��*ߘ���is��ŋF)3]"Ι�M]����8t^b�͊��7�B�~#n�@QY=�b7X��g-0=�idH��9��qQ9�6>��
G�k
q	�����D
vaH$����WnǬ4�Vy�c�=U��M�i���s�����53UV�����>|fG��z&��֨㶂��?F3�'w�(`Q<�2��Q�t��3 �z�>V㊁��j�!�T}��vR#��K�VŦ,L쌂2f2(Jix�J��2b�l:�h��+�#[���V�r�9��a/��2���R�aRN<�X������{#	A�/�c_E� �e����[aް"=�j�Z(Ep���X�j�aG�w�.�m��	��T�s�����l�0��q=1��,yŧ;Ѭ-=��%� ����sa���^��%�%\R�V+h&-v��HIuV��q�t������\�$`�$�/k`t�)�[�)��:�*)���.J2��eKm/m�� �c)��n��1l�~�x.��u�(��P��ۏ(��SW���m�z��T?�X < EA ZkJg⑄�%lto���<�IO��)>�a��Ե�ÖG�{�Q^���0[kE느����Yt��|��!��������dTK�z3��H<����Vz�K
^*L~��F *��f�_M�M���p��g��E��'�L����xu����#嬦��J~�U�(�z�ٹ�ͺ﷞���p���f������?��G;�;��;{���W�?�^�<�����[�K�g�Q;�$?�?{�r*k��Kp�):_ã7�i��Í����n��u���W$!��=݊V�V�.@O�8>��X��#˝�O��+��Y��8y����O�7��J���˷����T y:�u������?�I��\@�Y�?6��}�(>Љa@���~�\�m��s{Y�euDU�I7k�}�cՑq����M$hE�����S0@����k��X�Gt�ږü�z��$7�म��i�����qjɚ�Q��1a��"sf`@��kt�X���AΣ\���j���!�ҝT�tz�7�Op:���Ǧa��C�<Txo��C`/pTp�T*��X���pi��f7����H�6C9q�<���w<�1�q��8���m���
��#��Lz����z
�P���6P�����K�3��͡l�"��z-b<���UZ>�`+Gά�LC�鞕L\�_�{N�U�<�s�|�:�u:2�g|yʝSf��؁�V2�٩ǛS�"�<vW����T��V���3џ=0�������h*�����0�� ��� �� ����?����.�֓�ΰ�_"�#;�� �;���Z�O�:�V����Gn��K-H|dq䦥�#H��� ����[K�?�N�O�+�9��.�F ���&�\d�u�Fj��ER�Fz��c�?���o+)4�������}Ͻ�4|٭��h���k�� Q<���DҐ��Ke6��8`�lXi����At+�"G{��?�f�h�qUK6�I��/�3�����;�^�"$Ř�G��/_Sv���b{n�ө��B93�Cl�?�bc�R��9<��'�j��ʵw�n@y0��1qƪ�&�����?Զ�>�D�� �(J��	D�X��`w8��R�*a�5ΞOk
�s���Խ�?� �06�V\ϳ�U$q��nt7׭�򦮸�����}�SX�7~�J��k�#��z�ZK�V���Xe�F��s	9��^Eo5-��9�g�ʝ���+;�|���mJ*$'��a�:�� I�"r�\�j���I�4%�笆�Qһ|tI.2��ƻ��L��-FW(��2�y �$uͺ�q[�����,t%�E�tn�ff�>��v�}�k���v���)��"!�"/����
}~�!�7�T溷�H���_N'�OlS�/*ڮ�?F@VH��fQ�z��!��i��݉:	c��߯�<ha�tD'vS[�Æ�#${0�e`���̃��"Ak���8y�{��P�7n�|FsN|�!���ˣ��dyu�q��(a��j����yW��H��)٧�o���`qt�/(l���'( I����DhdC���*��b̃�}u����E0��3�r��#�Q$b)�0���@5�_���ρ=vJ~����������gl��C\�� f����e�B́�{[�+@[XY����,��^��>}��mT%e-d�Q+ =�fU}^o�c%v3�R~84���6 ZJ!r�_k�H�16pS2�1c?b���)�x����������z�$W�T��f�Ω*�\�}�V/�W����19����B��U�8k|%BLLV�-�W� ST�w�ηv+dAk��~��F�l���݈��-IϮ�����[9�W���t�O顽aT�G��b�5B����IW��H%�U�0u�1A��`��y�����(��*����U�Q�~�2�Ht_*%iC�e�4�� Ų<)m���h���'����d^�X��o�:/^�����㗖�4,���\�1�w���]q��p�'�y@���n&�oʞ��0���#�x!e4���$ts��c���!~�<'�ϓO�HdBi{cp���3��V�=8\=���Y�Rww����b�}����?��	'��?�m����ixۯ[�ά&��@?S�>�Ȩ�` �	��)C=�Ly�H�qfC��L��&�yW|Q�l0@�����븚t������'�$����,��nv���f�Q}�e�b���ȟmQP75rB�;:�F�|���Ӧ�MɖH�Y#k���%�����(hP�F��d����3� ��{���X ��'?[�Y��#<���x�(mVU�q��A��(<q{�Jtis�=DZ�{���	���Ř��>�y���?���i:�5��Xc�L�{\m��
eY\p��5�E�7�^����k���n<�����|�C�Pǲ���=؁JU��U����&�l!)խ�o�<�b�yG�4�yƏG��6g��ϷJ "X���I1;��s�I���t8>j��\Rt=G祟�����g���.D�c"2(YW���K'x�n�y�!#QW�A�U~�6�^:a�q����j��tܴ#��CԂ7�U��> ��Pi���\�4ȎԚM~���{rҲ�\ߕ��y����������B�ʇ��:�kS2K)V.�  q���f�����w��,�l��V2��r�����v����@�*����J��7C�.��
`�/��(BU�� �"KC�MZX^���8�0�mC��j����Hg0!'��#��8�����J1Z�
�U�0Z�o�����fU��>K��-	��}�if��K��բ�X�5P�ʸu�6�1t��#��`ۂ3��B�B�|
 _3ɮ��^#Ÿ#�Ѓ7P��`4����w�0I�Y�ʏѼ��Y�'�[�E��L*��W��P�e���0(�x.%�0Pn?�<9h�w;��E�?�P���� �GOMoo�d�><�?ŋ��}i���ߖ�H?/�WoY�ⴳg"�Á�o���G}�6�U���"��;x�_����h4�x��MP5�4E��˼���	�4�U��<�y�M���f���*�Zw��'y����O�W<蕝����9&e�☆�}�M�ń~-��Hˑ�-���Muo��a�(3Qd|���wq�����S����n&�I5�R�8�o�%#i����aP�v�ע4Xli�Q?g�1���rA��	Dr5��W�i��3m����v�J�/�Θ�`M4���� �C�x̵f���� s�V.~���ʊ�->>"Tf�L�Te$�e�|_\Ev�c�LK�CS���o�Z�p�{�����K"`w����q#��_�?�Ѕe�Wd}��y��$����9�ηs�/��w2�$xT�ߵ��_�8#R��Q� ��a����7���Ҵ_,��~R�B�P��������Dƛ.���D�D�(6����&��UN��q�wi�^�/Sv)�^���0.�����y�L�\K����C�U�}��FΗi*�ĕ!"���i;o嗂G	TԶ���Pɪ�!l�Q$V���ң��B���S�&�*D�G�%�;�$6�Ҧ�����n��n����X`�XgL�Q���@�C.*'=!��_e2g��2n��	���N�T2mm4�&- �" V����,��ȣ���eu�Np���G�̏e����L�,��"���ǪdWE.�]3y�a��ݳ���>�rO<��0�bx�������+z��`()w��������A]1����]����η�/rbSm28��h?CD�Fa�8b�w�7��|��Tי����r��O�r�?� d����4t�� v�ܝ����,S@b܏���MN\�9��Z��S�#;+r�i���=Z
�[��ظU��:Y��ߓ٥��ruW�n���u��_J�^��ڻ/�4����t>W|�ȼڋ2��l���?�_�����m�x��J]�oyh�����`8&���!������٨7 FERp�Ǎ{Z�{V��ɬ�>�*dX�UV�s51�ry���.�ZzҘ�蕘������	�䢮
��2T��=���X�uBpD1�h�L�n�D4���"�.Ef�|�:lHJU|���sA���u|G_��{���\ؑ ۇ��jԑ��]�}�R+�6��&�J�$�v&�g�:_��Y�9��$����+ F�aCWYM���zWtĚ̙��%�������v�_���g9�Mѐ<�ɞ��R�G��xpCR��M��#E\U��R�ܲ��Ŝco,f�4��eoX~�5��C}���U��wp٥��`�[Ꝑi��'x6��;� o��Aѷg6����f�X���ʇ��'!�ő�\��,,���]�r#�ܗ�ÏO�RGoG��-x�֧r���ńi��;Z���x(�&��YXuϓ�2M�|�' R|M�}��N6:5N��Dr���[K�����U�Q�ɂg	p\d��y����W��Z��w}8�'���l6��$�-�r5���{(��)�=���Qe���=�1'���o��y}��1_w��4�����U��zzJ$�Ը`V�G/�6�֚?�M��N�Q���YS[O)��a��gR�Ym`��:Gi��z��sN�)B
�|���;�-A򭋜���>�Zu/�n�-�,N�'!Ą�$�cU=%��Y���(G3�C�\�m�ŷ=	H�=&�*�DW4G*"�B���Lz1wf�d��ƍ�4�8x�0�c�2
V�ă�sk^q^-sn�����7�����t��|"�6	`�lij� �o�jOؤY|v�9Q|�g��U'�5��߽.S�)P$����n��M_V]_ޤ9��	]F�Oi��������GOx|�<\����$�O�g�ݭ[�n���+6wS������T?QZ�Q�j���7�{m״oW_�� {���9|��i��M���R�i�$e�%`[�7�G�
���AI�����q�"�WG�o[!cN�1�!mSw�l�>F�{����?�l���Q_�	|�'��ed-�"�ə��4%�,����Q���6��+�>�S���ɑ�Ь��k����$���Q�3�'vj�Ṙ7��-]��o~'��o��洕�Ҭ:�}��*9Jq�_��EP��_?c�X�e�\�Ojlu6���(p�F4�J�ÕS�R��J�t�4��v�΍�Khg6sLyu��:��.3��Y�	�M�cl��_���<�ݎ��F�S(\k��5��;����M��
��?�;*�_���j��/���.�>e�M���ɱ*X�m7K�eM%w���M\v��¹�P"jXx[������-��zA"��u/��*g.�
;k��<*��:�4�J̟�����S[�	KL �����
�9�����~�x�@#�D���)�K���7�F3���,�
��\�گ��f�咤���r��>cC��7XI�uD�~��q�s@�X�w̳)O��}ڤf�)�Ut6�լ��[��G�a�G��&���B���О�?���F�/E�Y�pI��y+�q��wǋ���gL߼�5ka�pv���ث�[�B��l���M޻��&�Ւe�p���L��C�>��!�]u��+�����Y�No�����R��8�]�K+�r6�{g���u��F~����-�;�&��s��;���[�
2-�̒d-1�������`8{(�O~N��`Fɶ�<@2�q-yb�m����U��S��<`�4����'��dr��]��rot�݇���|�;�t�e闿Moߛ��B@x��<�{����Z�]ӝ��9(��/�������T��3���*J79ugQ�W�L4���h��h�-��RW�<�=G>t�D��Js.�Y��T�W+���j�%��
��Z�:��_��2�NŐY[��c�����hoe�H؄}���F�l��J��g���x��	?��/�uQ��o
_�9�Y������]#�<�6�����S�>~�gb�!*��.ZM��&��ֆ>]�P0�sf"s�*��"O}�]Rɠ�2K�5�۹�k�y��x��@z7�ǈc������Nzд�K�ظ%��>;R26Y���i��d&N@���_8�:.�)�ߡ���	_��	���Av���6��ڍ*��w�bBFUу��̠�\!�.w�>���f�T/��u��!;�����Ե�ݾ&ăJah;O���>������sL����liK���	N
�$�m�}�i�Z±��J��r~t<��h�3?��8z����&{��y����O�x'�e �5�Rw���:��v�������[��C��z����ڇ�B�����/���RX$t;�w�e�S(n���ـC]�͐|�).�1,��&�5 һ�"��S�t L˟�P����R�xJ�	Bx�9ZF�,G�U�::̚|�l����_�Y W���9O�K���I��`O)�����	 �!Y��P>�C�)�6xck�+�}� R�{�.Wd�#�����M�B$(:��[�׿�ZQ���M���+��bq�wu�������F��dr���Sĥ�C��z�p� eni�L�n�g��z�$ޱ[5�4��.�H�\��	&y_{�����"	����C�j�����؊�7>}=	eI[\s��j��9o�ֳ��c�:�����G�=ėz�7G�9���
Ƨy �a�hK팱|��4*װ��Az���۸>�g�H�Am�H�;��P�?�2
I�p�n�����#�?�ݑ�6����<���Fɲ����=8^W��_޸[���hª�-VB$������? �)j��eH�b��L�G|J�9���c)����"�%{}Dn��2y��yӬk�y��]
]��q��=�H͍��u4�k��W �1�c��L��0;��oj�!Y�Ö����h�Bh%�N���QdJ��)���R<G�eKf1Ub�(���G���W�<��Y��8M������r �~#�jV���.4�W��h�髓�"@�$�x��M��9����7�R-�&\-�Fk�F`��	��(�撕n�aN$7��Z�H�w�`��� o�f�}���vv��f6
�l��!<|޷]vV��q�K_.,���.0��&�>���Rw�"�;X������f���(>#3�;i��繣�8�|e��:Њ�aw얹T1H�s��m�WW$��:L͗j�k�wi�I�B��d�1�f��koۯq� ��F�Y\-ӞM���o��Hq@$��ϝ�ӷ���c;~��유"¤~�'��&�^?e�.�q;F��Dt@��uy��X���ȭ�/o8u���r�����^�߾�StߍCA���ׇ�I���4���r3�d��wa�-��0�T��_rW}���L������@�J��jG��w�:��U�Sq��f t0�p� 2�~0��u����M��!?\�"�Ԥ�4��߃U�SW)�D!U����K�g&���t���߭s<γƥ��\�����L2=�֘X��9���o9��_�cw���v����^�����,������H�ʠ<5ݺ؛ڢ�<�ˎq����D����ھ��5; jk������wS����̪c/�Ev�V�ĥ���&cO�⒫=��.q6�������r��0˱��+���_1���Z&�C?LH�_@#B	ò\F�,�
�o(���p2��f!DÐ��^�`e����� �1�Uv2ɋ2�����b�v�<S��'Z��v�����,/��>L{��^�2)0����v���3o[蕋_���i`������m�xs��|�>e��̿����x��:��$W��d�����֠�~�%	λxC�Ɨ�"���m�"	�g��mr��@�{jH�2�@#�m�zL|+�8.�`F_�ʔ}M ��4|���Q`�����[��]+^q'ƦiWO⌣�_ef�so-��jf�:U*(s��9>~�AP��Ln��n�8%a^Q�RL5��e���I�9o�e���j�I�*��dӞ4'9�">�w@�0e$7O����j[�j_�s�em>l�B�}����l�,��_�M�N"ŜL+��q4��R�ԓ`�增t��Q�>��� ��%��[$�d���{Jw����%��.��"��*aW9	{��MԎD~X�T\�_�Tu'��3�r�ֿ}޽��&+ts]��	t���%�p�w��1\�>����m9�c�":�����	���̤e�xi�Fa����riMٸ�����XH�K��K���
^�O9ULd�Z&��W�)�~�p��[Q��
�~#�*��rm���������;m>k�ޖ�9:��^4��[����u�\��-ʁf���P0�T��?@�vQ��m�E��d&`��`���ӕ.�	�KJ���1=5���%J0�+�N�k��x�$ʲ�:�~�Ć�8����lPJ�[km�Xp�dS���]��d��J(��ɢ��{�4O���$ݞ�>Y⊀gN�����Սa]Ah�ʍ�1k��4Y7~B��H�$�m<�;��F`���E�#�	����2��U�t��;n��<T����+��x4�9���M+�@M�A��A��T��'s������*��/	�-Ci��M� ���y���X�]����^ϻuz����֏b���E?f0��6�_�����F��Qz������݋�݅Vr�G�qA�ʶ��@5A�K{-�O�F���M�'_Q3k,pp\��ڂ��u
C2��3w�pqU�%�Ûd;��W��ck���0׏�~�i�<T�4�4_���*�`R�TƉ�k�G���e�ŗM�ɜ�5����J���غ�}��HI95c'�'��T�=O�C�Y�{�%����N��V�5�,kG&���1�=�aRߋ"�]�?X;�|>o�丏O�d�x�V�?43f�x���N��f
VВ��ã'���]����[HU��K��6&a�DZn�Ax��A�9 oh��,����K~��H�Gq�m�<�I���l��Y�t��rg�#?�cqC�Wrl���hFdr>۽Nn��%`
�M�x��MK$N�t2���+_�,o���Ldt�w�T��H3��;��u}�U����C�>���	'Ӫ.軦�er�}3������$��C��s�;�ϭG�L/��]��}êz��o�u�v[~үM�0��؃@Lm|ҡ��_�q���'�,�V4U��B�p��w�W�V�\�)h�RqK�z��S�q⠯��`�?�s���/u��-<}+s���2��Y�9!{S	a/�!�f�����J��VU��t�Cy��-T��:$f��<LN�k����l���v9�����%v�{�8NEӍ�U�D<K{��K(�R�+�����T�x-b��l��6�̼�3W��V�Le�����Y��qo���e�s<���iYث�����D���̇�&��y���2��Z��p��X����t�wu���Ub%&RGz���D���9Grh�����di��x��:�������6L_nRy�i/39NLj �*�C�Y-q
�H�.�)識?�e��&ѯRݡ��v�~��wwa�R����T��L�D!i�����.�1�=�E�+yN-͞!TL�)^��d#v��=[�n�d+R��c�m��vm2W�`�G<�^H�]��V��@�L��ܺ�X�t=��v-�\�p�1!*����7����\�xp��2B>(��7�w?UCH����Ѻ��*>N�ui�C�EG��<���~ۢ+}��
&��xV1�^�a��p�#r�\9.��*j�y��t&��g��=v?~��ZQZh�[Խ@���K��j����'��rg����2I9����m��x�3�#ek[,NӐ�2�/��]�Hh��Ud�pC�����E-����"�S:�.Ͷc{����F�VÇ5#�Q��M��昈�2VUx~�b <�<$_��r[c2�khz���W���T�95�g� ØKC��{ؙ��'�o�O�P@}y{5�U�L�u������𯸉K���068�J� ��񻙊ncF��Q�����^֝X�ȟ�~������[n���W �V����G�բ(�����	��e�
���]���hp<�UM��0���p��(z��?#e���I�rص8/����ˆ=�!)?��0�g8��ʽ�\%h�@A��șZ��`����ѩ�H��V!g��da�W���RJ<lJ�e��|I�ܨ�9@�ѫ��qƕ�J:�4���N�:=z,�#D<y/�A�1$�0�%���"�y��@
l�l{B���m�_utA�'�\b��z1�*�$L��XZ��yz��O�6K�a��e2��D�?W���ǯ�޺�jx�%I7@����^:	��}~4��^՛�%k�eB����M9�u�� �-,/H�bh_j~.����S�-�Ixf�Λ:�0R�0�VC���ע�Q���6�fʅ�����%���Z¤��1!};�B;Y0|�Teu ��(-�/>X
�}|��Q?�'֏�>������B��r�|� �o�;Z�6�􎯐,�pr�x�!���3��֞�ƏE;�����(WJ�W��@%)K�#?~._I��\�\E�4���U�*G�E-w;ON��5�l�*Xބ��N�}�M���v�B��}�ُ'Bk��{����w$�u0�h_��PA�3�;��3i���-���T$b���?n��:+:Q��j���g����p�Л��٣0԰���뜾	}�}���9E��l����_�i�Ɏ*��=n�t7=�w4���nT��4D��q�
��JH�	��Uuqc�Q �b�Z-�����9Z��`�u}�lg�'9]�M�u����	x捯����sĭ켳{v�Y�+�ĳ�q^H?+�����4������;'����Vլ�՝9�L��]
s_��s<�#im╌b[%�u�H��^��8�(g�y��h<V��˔�uW�����w̨��|x|�9D_��)�� E�\���[
����"^�f�z՚�[���{3Y��7q�C��bX�o���0�8�T�[��tk��z?�ͯ���U�U�g��
����3�v���o��Hv�ʐ��RtS�rv~n6��ܳ�3�� I_���78l#�j�Yg �ğ/#�m����ĸ�>�g�Ix���z�����/m��1��T�CH��s�k��<|Ia~��mb]����m��D���涓h�� g�W�H��,�%����J��@��Z'��>��k��h��>���jj�M!�W���-Ĳ�a���r���g8r���
T3��8�pQ*W�NZ�n���,�)|�0�z3���l��u��2@�N/M���h��c>9}�'nzN:>,m6��a�ſ\O�
.gȿa#���m��t5���G٘���t�#��e��r.jo�_�C�?����H�r-6�Wi+D���ߋ��>�h�_'*��i��}���Bp�A62Q�#���<x�śa�����1���ɚ .E+�Ͽ(�o���"��&š7���������)?�؅�G��h���ݐ�D�}]QG��-���ތh�vO΄%�3�\�|����S��|#HQ*������	r�,;T��~��]�LgP���{NR^fbr�ꉼE�󙿁#�г�!c������D�f���g˦��?��g;�@*��g�b��˯ע6�`���U�'[�0���x��Y��-���dJ+���}�A�{BWsa�]��x<�m$�Z��h��H�%�셅m$�^  l�Z��<�i5�����z��
_46���!oYB:*�E2�b5�8�1�1�ʄ�>�L��]���+E��υl垹D�_ޜ��Z�)9}�Dc|��U�at�>kR�ґv&�V��	m�����ٸ%���á�&O�o�?FI��k�5L�lxfq��A-/8�2~5}ڵ�C��F���sxI�4�!�gW�&@�3�<�)ϸL�]�J^+3\�l����%��J��*Ե.��8�� �aGRr6���0ou�<N�Jq�Z�}m]��9���K¤X.(9L-"�w��11b�Eht���=����*.�EǼ�]J5W�)��d��De׭�2��I	!��m��x~-�W���\1�5�n���0R���[�z��w��>����Et$����|T�E�B4P�0 h7����51J�����>+Z���2�[rS���|�2�*NրɊ˼1P��=��Tv���DppXZq���2i�O:p�~]tzBC`b�Q[8"��Б����~�w�wλ��)���?.���	�ٯLG�ʏl��I��� FU�ԟ �k��
x�怜&�2zA�����te����\�Q��X�jksP:��;9�2<b��n�--S��G�N=P�K2ޔ�^�ڴ��3�g2J��&����OJ�k��H�:\���|9tc0geP;?
v DG�:7B۬ņ#L��h�os��0$�*.�! b�!㲴�G�x׀�r8�A�xgׯ�]IMl7�溡��!i罜�ӧ1��J��k����Q/��l�P`��%j�t�my12��>:��wB���<g~AD�ȇW�8���SB�����R[ڗ��{�ea�s���d�]�?��g��^[�����	�Bn?��{ɠ�"�êۺ��S_����:�����2300?f�����捔t����u���B�~�'�7�C
sc���n���4I�+�x�`��.�3�nh����Y���}8@f� qf��v�2��%�x�t�u�$Z�FyqDM�:V��}�!�BN�7�&<ȸU��!f�����,ֽTA����M��[V���}���9���L��ߝ���y�r��El>����n��jh~�]]]���i�a���nY�0�w������3չ�Q�O)ka�0Gm����O��چ��P`�SU`�半b<S����y�]+K��)I/w�e{�~Y�Q�@�Fҭ�=���{Rz}3��ދ+/l�����3�E�Z�lj��!���HN<k�g^�և� }7�Jҝ��AҬM<N�^�vfa<|�<^vr.�}g�9f�#h�RQmU��4� W���{����9n��#|洿�ӗW3kj.چ��,V&�J���EgV��F
�ʉ����ؔC2K����+����]u�A�V�_��[y�]�\pR����R`����x=!� *���G銜H�! )����*{�r>%7���N$Y�}�#n ǁ݈H~��U�a�~C-ޚ��{�LDe}�~�Q�A���Lh�G�~�;U��i�.8:��Q{��|��@,�L{zE]p��O��{�c:-ᯀB.p�L+�p��Ii�O���QK^��0����ˊ~�*�Xυ�Y�ו(!���@�t#(X�{#+k�Ƴ�>�'�-�_�{���?"����`���P��pS(�������a�YjԬ���l,V��UC3�u�Y�E٨��dEZ�WW�I�m'���I_�SuNd�����筵����jW�-�a4����/y��r��LlQ?��ҩNM��⅀�Sb��G3�N ec�ɡO߭��e�����Q�/��Y1�7�DZNv|6��}z� �6L�R�lJ&�ҙ�V�0v3/�Z��� ��� vm&�:�6���P�+�b�G0ն�1�	��5ș��r��u�s`O��JÀ���C�8^��5�;ވ���/�m����1��r)��u�a�Q�U��P�׫Jp������A]rD]#k�`��Xe�L�VD�H�Ԧ]��4��*��տ
]�=&P�x�W��pbz��箘���}���8�؈�#]M}�p��=���vq�q��	W�F���(��$9b��PS�Gz��?��$fQ�c����N?_gA2u���%�>-0�S�P��6���s;VQ��t�_r�H)d �����?Aa�t����~� ��߰���D��d����J�[ D���ױ���j4�x1M����U�<du���W��%JS4ť�������Zj��e�njBnp2P���nP�gIiT��(�'`��;��sқC'MFUl:EB�Cޡ,%�YَL����A�Z�ӅNy��C����#w���n�����K�{7���'W�^xԶL�F{I	��� ��>d a���y:s�d�M�L�R���W�^�7IFc�e�ڢ҆gS9R��=$�w�����F���~�P\b�h����A{�'�LĽ�������c�_HH����R�����+?Tl<%�^й=�,�>�sMӔ2q�)l�\���FD�@P���(�>sY#��s�T(�8DC�,������� ]��d��A.ŉ�p۸O��ooo髢1����i�җ7,�4{�E��5Lî��zisP-����3��yEv~v�٠�:�8[;UCqւ޲��v�MB���i }�g������hK���7g��*��ϻ�B�5�?חNI���_*jF:B����08��(�\���d�`�{�z{��L�^�zeSK���.p���TVE�d䞋*���?OfIn�`/e������ �?�HK��7��T#}�R�Fv�@?NrsB��)�5߇g������@Dh|=ݾQ�y���0Q�+ɣX��Ƕn���[���䭕�)8<C��9���/)>�-=��K�x�>��MD"�X ���	y׮���t\�.���z�8q�����@�B(rB�x�3R�bc�.W��M����w$O	��+n2癬'��Ql��#%2��������[ ���N�iT����.�[<��g�Į�%�K2pJ0�D��-�u�B��N`�<��}�pjTN<���#Z�Q��^a���(��l��|�E��E���ñ�(�o����&u�N����Ĳ�f�1lFJ �@b�8?P�M���*%�il����SX�e Y'�<�Eڋ�[�%ɳ���<929�u(����y��52l�:�$rH����U�� �3��5-?>�r�iA�<�=��	R�@��PB>Ņ���-���eFSw���������6���K��fD�T!z�����0풖�#�b����+�Ǉ
���YQ�}���SWH�.E�'NL�����T(K�Ű��^K����c��9�~���H���N�~L�l�r�zx-�ϯ���63c��If,��џψ"�ԭ�*��8rf��[�,��I��W���-�K%&
!���.�����2N̕�(��?#���[ɲ�(�v�� �@#�h6��"�Yb�Im�.fD������b4@�0u�ӨT����rL��H� �#he���XO.&�&M����9����[�4@8t�o"R&5"ށʼ�
*����&L�'��󘽊	��S��\���pom���R8�%�����dْ���Z&�fD������h��.x�D�iV�S;*2��P�-�%&ujc ��̄��8���zC�K�w-:�b;oo�0���t!g�L�E�\}Cou�ļ����f�p ���k��$u�D��-#�<k8\?�ujI�>�~�C��N ��#��.v�*+�ȏ0�,��WAF� _R�v�G�e/p)����W#������}u�X(/l�OO�Q�I��K/�F�@�s��A��"�����'�:�|�w��A�n(g��Gq��qj-e��0.h�3u��8��ngTdax�$�"y��ǿ���w��ԓ�.�����XK2K����o�'ㆶ�!Ð�8�Y.Ѻ���L�(D�Y��q�v#��@
34H��A@��7mҧO�(�ڙ��)A0���1l��Q&;Ԛ�Dĕn��BE��C� Y�aE�nn�	Y
�sA��ż�f��&WEO�b��(�S5M�����V���Fv&R7�v��Q�$Ԃ��>!�g�i��@���"f���B7�9)����<�a.4�.T@D��E��ʓXm�B"A�f6�!c�+�f��T"���N�`P!*2h�K��Ɂ����������2͸
�O�*&`U��ʼ�T�z��^0�:й��%�-�����y|��0��?\ty���4h$�s�>���}3�c��d}�?�.sҡɮ��R_�O����'�m� �n�?g��9C~�9�l�]Ϛ�E����u��+	6H����C��q]�X�]119��
P.ShDǌ��D�7�B	0nҟE�BtJ��x����ۅ��ﮊ��q�B���3{~x�W�71�`� dC7��Br`�������^q�ȸQ�����0�Iߙ�o�L1���\�8�dXz-�r	� �V�������.�`Q�:���� �����F@I C>��0$e�;!B"vRbL!�J�-��E��9pa#�C��X��))V�VD���"��ټ�:}���CQ<����y2�� �ie����d$$�KH.��,��8(�����!kl�G�n,Ӵ��s��6�Qt�F�#,*�*|XC��P$b!�ΣF9ܪ&	�6�9Jb��	O��W}��/���u_��A�^<��4��7>�gHǎTz|��4W�Q�p@$�)���H!j��a�Cq�i�Ei��f*!�a����h���|~?���·�<���2���7vv��.���jyI=!�Ɂ��.�L�����i,����uL�m��̟�����<*y��)���]@�|��gU0�m?9H����y1�RD�|�a`Hu��ϔ�0pah�u=b�I���_f���Gݙ��#/�8��(/(� � 7�NӀ�Ϧ�0�����S��,�R%(O�?���pr���p��l�R�5]��B6J�w%�H�։X��<G�Dä7*�{�j"�3a%�b���6!f<b��IRQ5�ik1y�*x7�C��
��r�\�01*,�!��o��EQ�C6i,*$���q�(� ��t �D ��
E)%�D �m�Ӯ�9)�(\�GT��&�7'W�M���85�(�B� ����f���v#v����elሦ�	�t1�0���G���1W�o����l�@J��������`y�ᒹG�+�1S ��i�	1���!(,��X����~q�PG�oD�?)�7�Y����r	�~���S��0��c�� ��ȍ�_���/v}=VgY,ɾz��6}0��F|FEvvd�9�9$6�I�L5u3�A����4�R �ew�I�А����� �� Mxe>���cq�k��;�Ƹɏ  ~A��E�H����#SBϗ/�4�bK�H�Y�.t��C��&��č⼸�yc�;S�%�W6��q̐�S��a<�7H�a!�4���������{>󆢀]����gF��
H5��X�0��b:���y+a5�&����p
�@�� +��Nǘ!��I ��Wa	�mHd��!�de�,"���H�s$=��� �&̠�F���y��Ae��;��!��+@$ؐ(���JlD!4#�3SY)*IrFN�5$�LAv��(G9DM-YS1䣒@AvyG-����H$ks� ��1
�A� _w�����-׃�x������n�`��a��Ic��c�ͥ�8@~xd��d����H8D�D~_Z1��������? ï��_���1���-{_��K0~/�̱c_}ØAS?˴�o����"�ɐ12D:GX����!%�K��Y�f}ܺ� ���|+�@ �,�	�I0��Tө$`�<f�D���������p�.\Ee$�qw,cV"��We�@�%
h	�ry�LU�����K�?8�����?����.)ͳ� �&hyk��ej��.*<A�m>��8x�Es6�Qu��p�6�w�؏���<�6P����8�jL& D��NFH0��J���Q7dR�p�l9�$�Ā�hh�Ĭ��Z�#M5ႁ-�\�y.[x���ܬ����G�F$jow���F�JI��q%��1a%e'��}�C!�7�����ƅ�U12R��Lz�,"����1D�z�r9m#[I��2]�w� {\����T�1)�ĭ)�G��弆~S���Os8A�����ȑ����^�1ƹ����q�W���*�	���r���v��'8-+O�����t࿟��Dc?<F(��-�p�� �mƬ/"�s�5������4�D�J��ND��8�Z�}mW-Z�B�@|~s�H��8���2�	��̀�"���F!*oOd�n�� V�22`���d�ց��A�"���2���}3ED������r��C�A��b%1(����$�QL -|C�!H	|'{&��ntI��L��&D��R߳���8��/��'%\�>X�N$+�,����1B>�:,��i훎Y�3��௉��U�a�1��s���D�U�<��Rk���4�&�f@�Sڲ�)�0C/���jJ� AI& ȏF�r�҈h�"%0���ndm(�#����k6�$D�NJ��>�	�}�l�J|�B&pĭ��3��d�|�߭\��X�M����*Cde�+�
ed ���Û.u�%�h'<�q*+���Ē|aw�-Z~ x�g�?Y/�r<�P�|B��5 ��tZ�T��l"$>�p��1��(��Ⱦ�?8#�K�N<��k�ɋ�;�������t��f������h/����~���a�ȂJ&�J}0�J�aI��q��)��o|a$�՟.���E�|��w�G
�%�czL���Qɖ���
�r$�*�^P��N�cx��W�x��`j���'��bY�J��;�&� �����d�����B��DN���4��<��W�cs�(@��]'�����c;� 9���IH�O�A���EȞ��&��N>��aT�LU���x<��8��6���'�?�`�9>r�� A�B��*༭�3��O8�Ϳ7��Ϙ}���d`���߱LTMP���`G�-)���U��',����Hr'a �����a���p�$��������� ��5�C�ۡ���>ANB )�b9�)�T0�
d��2�JaDE~!���NM��������
<�B�1�%��6 @�a�T܄��U��|d�u����\�*�J�G2t`�PJ<z��'���_�Y2�eN�u�o������U�t&>��G�Ů ��;����������EdK�p��+a�ײ=�<9Ӹ��Q� �,ށA�Q�Zz���Z�i��(��_�rgF�H���ϙL�S����� ��:�0:���%a�C���·h��14���dNbI��.s�9nO�?��� #>.�$�������$�A���Ci��<~s���ilOE9�3�	R��cd���D��By���"�<ɳ�, ��`�[?�� �W��ٝ�:8;��OQ��;.A����� �]1*��pNV}�������&xZU�:4�+����2U -E�`+x�\�����`��q�VW��c_c� ����N(Qc�������Ba��	W&$�����'�	����G�� Ư��D ��}Q���a���Z5̃X��k�O(N�D����H���M�,3@�\��J���P.��QӉ��c�k+ғ��kS�YT��moW�%�zLJ�KC� �!Udq�5!'XMc�$DÒ�l)j�K
�t���!�2M����HF�� bi�2;�W��R��ń���!���#�`�of�����sK�N��|��������	���p��H���E���L3��_�5>�xe����܄����䗌fy�H���PW�k�.�a�������lBw|�=d +R���S�?���Sx����͜V|� $Iӑ����|#YO拄�>��d��TW�D�U���A6BG�g�gD��������+��~T#�i;'���3���Li�d�h�)*4��1<Sɹ2D�O��`m��a�ĪnOQ'6XXn,&V�NM�^������ɕ�}��θ�2Iѱ'�Z'4�#�U�?VS,t�`sxo�Z�^��8��V�,�_L�B0Dn���I� �D�9�gl��&m�/��fH��4�؎�2��!���:�6a���^Fه[g�}��f@�@K�z����xȗ�7���I- �0,�2iȿ>ĺ�l$���"�dy�:��\��hx���2�=��_�k"d�����Bm~t��0m�o�Vp�RU"�2��َ�0/-��HK$e��%P�H�}��"��D��(y�u�ɾ�\�[)�:���� �DA�A��{P��%\݋��&=_�	Q�T�_�j��`��^<���vu�bZ��Ä?�y����(���������A��팥�&�� 6�Mt'��~`Z�ATʥo��S>��L_y���k�\j)C��dWʆW���8��"�.x	!j��Ǿj?41�e�]@��������><�G%(@|d�1�wz� #�?��ñp�y2@�`���a�Q�v�����F��+��1���� �wZ�-�� �\ǀ��+��C��Q��VX%D˂�Q)��i�u��O��6]����da"RqH��<&y؉�����>@�t�E�K� (��uX�L`�sn���E�b( F`4a�eۇ�"6+ҊU���7�KK���(;cͅ�<<�V�.SX懂����n�t@j&y��=���.
j#�πe���YTu��M?����H�5V@)OsS�31��+K=���d��g��"堌h,o'�U��� h��(�$��Į^�p8���I�.��b��HT��o$��	�1�{m��c�Ʊ�K�Ϸy���(�$�\ó�ؑ������<�����[e5���A�c��BP����9la���	��%8 f�����"��0�q��l%���A:M�cl��k�?k��Z=O��~.O�N:����F8�
� � � ���a�˝{fH���S��Ko�{���ѹ� ����_��A2�*�K�FGv9[P�w'��"<�2L��p;:���-@6��K�Y^��I��O$Y"��/q�ʡB��I��1��������IŧOqRy��v"LF��K��O���#N]d>I���s�'�Ž"m/쎧�ę��"���;�\��L�y2u"�!Q�]��B�$�#:r���5��`~��� b78Y��]�eH�����;VԢy��dD =�[�dt!��[�%w� �v�q�wl}�vzA��JF2�1|48>����H-��8��y':�Ev�L��0�ľpP�@i���nri�=�r(�,N]��I"���i&&IZ�DB�A�&���t(J��/��ͫ���j'"bp�Ѽ]�zq�4=��4l�<����tB����2�����a�VL 	:�<�?S"��ᑓ��W �D�L'����;��D8��^�$�:�}���nۀ�y[�8!DW�!�b��?L���/����G\�#��3X:��N3���o�W�.�mOO�q�v4�� �|z6{$^8���_n���~|C�_��dz%5c�� Tl�$y��C�qy6;��'�C�$˙�AU/����v/�"5�Q��C��>͙VÓ�mO.Lz%l�R�x]�d��q$�3t��2�nW~�&'Q��{�	%ԋ�l�|���dy�9�jv�N�q�(��I"�a�B�ʖ�4$�f;D)�U���Y ��l�`/p#�'مA��Q�>/�6����t�!/Y�(�a�Щ9�`���*y�c�8�*
��r��<���*IJ�}^�@!@�d[�c�5�
^
H�j�$HD|��n0D�
y$�E9��⸁"d#�Ѥ,�Z�A6�by�-��
���Ĳ1��J"�͝�'r��:R�z/�屖A���NT`nI�,�����QN�4�Uϩzb����lOl�d�=� շ�N�:��|FD��_\ &Ծ*?X����5?Q��O��a��?s98B>�LUT���w0}\�{96����s)�@�2^N���1�n?�G�o'��o�g�Y;I߯umq�����x�y���s��}��>X9�~��;/����h9Pɖ�&������O�0���9�����Ϭ��w� 1�����B�Q�$��dg3�����B��T/!��,#6;�9������-IR.�1Ӑ�u+��-�\�(x݇�<������&} �"~��S1�<R_��å�HՌ|ۄ*%��9�2g��p�G��&@"f��̨�Ã�@�����T�ˉT�:Xta@���*x�ȔhiՄ�M9��ZL�Mߍ�/M�y��<"�����!�X)s���g���˾#�S�,w���6�3�V��K0D���:Ƙ�{���xG�  �
ʴ%�Ot�_�r�./4��Ĝ��	��p��Tn͘9u�Av]X�
q;7FnR����2F�dƭ% 5\H��F+M�er��	
^��<o��}���P�+Kg�1/A����ĢC�@�*���B*yb'Q�' ��n$�Z����}k%?�dS�������Q����r�}��`W˒un��t�ۣt�2�?���2؝�m��|�:8�9~�'�?����F��A�� ������a���ɿ���<ᓈ� ���a�1��%�:%F�0�1��8Uw!���w�w�G����y�w֡ĝ���`��G���w!#eVB^r�3����:-X���trvE��)~2���y����I}Gb?a��B���A�),�n%�����,B���?Le�*5�^Bf�	j���S_|��!�w��+y:� �{�"�l�AɊ��br���ɕ�� �+i9'(��9� އ-��X,O��:+L�2������g0���D����x���C�� \AB�@vF�w�1,^�ic8����1R�*hC���p�}�Ƣ4W��K�N"�1cu/Aˍ't�K0���``म 5��Ή���7�Mt��L�����L���$\���!7i����~2R��C����xɄ'q�;e ���^;�Ha��ޟ�MxƆ(�ȀŔm��"E>������nP���[�?,������7��I�J�N  ��y��{���yh�ID��D� :��TSDZye�h�HP�}Lq���z���}�P	�0S�댿\Оt�ǃ	�Tc����aσ?��7�Ϯ�D�V ��bZ7l%�Pxы�k}{������u���8,N/�w�*��epb�����;� >�|!T��w�Od2R��I�3�7^����+cq�sцv��UH�=�2,���7.1!���s��C,��yTb�`��i�f���'��P���ȉ��m�$���a("֣��uw��GZ�Kr�m�.�l Ө�� EN@��c�h��������Ò�5jS%���g���F6��0 گ��� �C�te��o+�����(�F�/U�!��L[��~V�O I��ʄIDF��E��0������jF�1�9nx�A>)��N��fl��e��:#����m���VR� �� �)/4����!t�^�_Y8�"ڛcp���>њ��#�Q�rN;1&Q �{����w�'�)���+!������7�@��yr��'Ì�L���#�%�n����z`s�Z�̇f�r�B�p�6=K��� wrϦ��HR����A󜩻�Lx��O��~�`+�����9~k�?Y���(�P	�`�-�8EG��`������'��������/��Gl�!��y~q y~�Л�H������Y"�qZ��'ؑ>��m�|�9'�\g��Zx~�aSr.'��c�)Ou��'���7������k�Y��+O��pzd�bN��Ewx�u��< ��DP2��ئ3t&�x�_l[�jY�o�"5!m(����Ef�*��r�L~L��gGeCɎ�,��#A/,s�ՋzS�s��W- c_�&"$�OЗ6�;>ï]7�(*���/�"!�\�,:kEi��Ő�V�Z���d�H2:�ˮ�đ-ޗ���Vp?�~�pή�m�&(�����.G���A�T �+�a2�O�B���s��NE�~��>5�_�~L�������)�u�%��9;X�` Qo�4r$�qP������Ϊ�>�#�
u��D�G�[G9:�� ��T����`遠�8g�_�!�������9��O��2sn0&�$'\3�`=2W��Wao��c�Ǹ�=z�;�6���> +��
zLvhxp{�<�x���P� Ī���x�|a��$���6��2�zq��GO�ѐaD�]��O=N:]	� ��[e���O��&�`��(yq'陝"���3����F�_��D^�>�2z5c3-��� ��ȋU�<�����Fhg����,S�;4~��$�H�>���
�A����hW%�T�T}���a��;���r�4���FB|�=\�.B��d��-Aܭ3�m5N�h	ds.3 $�tz�=�U�J'j�@k����I�8 �jk���ɟ��Q��9�i��_�C�St×��LpU�� � �a`�Yz�1��~���*W�.�1Ʈp@'��^�μ�l� M����F\Ѧc5�+����)T��2�x�`U#�`�Y�^V�/�T2�U��Qo�2F��9s����4����=&+�t<g9� ޯ&�c�!Gj��_g*���Qڕ�Lx� �a��D��+y���ӑ3]?�	���⏢�\���i� ����<!.Q��r�,�d�L��C)�x,�o.")U���8Bd!�W=�X̄�5��G�ee�^Y|J?8���%�Ǹ�Ȉ�r�'8= �ki+�� 0�K�*o�9��	3��*P�8��8�&U�V��II��Tڗ�O%�r<�8ӷd�XjZ�g�K�*.�ѿ����2i�oǼ*�ӈ@�r�1���,��(�V����A�
O���F0��GI��@�w���! A�!���A�ou2��\�����W�"V	���#q"��Z���A��(ȅ���ub��DT�w�3Ӄ�B��4�y|��Z�Ve'o��hܼ{ŉ�{�rh����=�vM�4���Wa}�BK�![�q���d���禬W[}L�c���E$W��.C����?�q����	f:�� ��tdA�K���'��:�DS�4�D�NQY�}�����+� ����P�C&���g�<���Y!��'�<��i��⼃�a�{���?؏� cU��T�P���i�����~���2����N����a��  � �/�)6;IW�W��@mf���4����T��A�4�x���,L!a`/c�\l��޼��0��>�l�}���*�h�1���q��H2H6��nw��@n�#	i$�F����9"�|�يC �!�{B�)���w��Ơ����'I�)�LQ�{��8�6	,K	I���L>K$!��N�e㽰6��-E!c�s�����H�W�=dH�������#���Q�!�B�d�}���IY}�t
���cW�IEu�ؖ�^�!����y�qQy ��N	�f�� E�u���� ����ܾ�����5^�y���n��+q��š�agݖESE������~�0y�q`�:Π��"��}�N��`�	#�A�g��s�&q�k�8��m��� � ��˖�>�=b�mC�,ެm����� �d�e/i���Rw����|aPC���&��+���?�4�q��X����pT��k�c�{k�ᨽ˛���i�+�`H��n��wm� ��G,{W�.!Q�%�,�$G�dǠH�����������F��J�q<�L�G�8��<��I˕c[������>��.^k��-O���c��r�����JqK�3�%O���C�$O�p� ,D�d���\H��;1�YB�O��c�����;�o�#)	����'��p�)v�B
���M������q0p.� ���(��lk���I$��}���BR��H6�'��81YhJ��$l4I�nh묹�b"�a�R�.��"��JV�IL��,������baBj��t�pD}	� �:$��cAОd�ĕ���'QKLoP�|������~2�7��\��~0�������0D��N>�GZ�iT2�����aU�+�=�au4K�W%"kc��<aᐨ�xL-� LxN���hf=�~�1F��[w ��-�F>�i���`��ݜ~1%��~�r� �����!|a�ʼB�C_�������OL�H�r�BT��+.�������0�k׽��xc��^2q]?���~�a&"VN�K����C-sH���1B�`��-����*�u�� E>\-�58���0�~��eD$��Gz
r<��Q�W����N���&�~u���z�&����ra �pby�M&�8�T��&��BT���xaQ;��\��u0��<A�����FJ��q��QDLz+D��w �k
���|n���1 ccd�D,�K�u��X	 QN�Yq�P`#c�Z�����a!�q��I勋&  � i2@���'��
o�v�Me�*�C"�}�E�pjCMm��Ɏ{�����6�~+����y��k�ވ��ʣ�����%�p�~�IEmw��aE���%T��ě��u�P" ��`%���y&��k�#�r�Xp:Z;�KF��VP�v��r��d�"I�!l�D��ɦ��_�K��Ns�A�`��]��,B�t<�\vC���������h��4�E���	���� �� �C�� �s��s�{��`^8w�͢��c$y끵~/��it��~������Z։~3f��A�b�������� �>\���*�7��k?&� B�8X�'��?g���P��VB,��}q�	Udx�����3r�KH�c�?��	#�k5\�ӂn���q�
}=���n��>���%�b��I��)|��B3�r,��f|��Yc���5�-���ˤsi^�@:��aI�xm�Ds��#`��$����bT)/Scd���R[R�:b� o {91��:�� H(��8mQ�EF����Sk�^Gz��6d��b{/N��A�48��^\�|�B-�8�%���N����q�� ����nw��9sA� 
Rh����!�yP�A��Ĉ�h�`�@9�Ȁ<�|�mb/�,
�Z�eQ,nX�(����}9�x��ѓ�Y<��0�h���ɒX������?�Ⱥ_����F�|^q��3N�?*S	}M}��� @'��CO�}�����"H�䧃R=�{Z-@�AK��EG͘BiL{���O���TR�Ez��7��N��k�-TS��6����z��CZO�!�Ł|eA*�Qg�`BsW��s���J 0y���cJ祿 �� �S,O֜�>�őd�<�g�n��m"cI��r�J�PzȆ' q±P����q(�� �������l;[���fἱVE� ��D�j��PD���d<	%�}������7]�����[�������[Ɇ�b�o�x�ʙ7�#��Dd�_��� g��}p����NAw�t�G�Ƚg?�&W���ϓ*�i�>��aQ"�0�ёʒ�x0�8Q�0�D�+8�1|�6L��?�V����H���P갃�6��O�_���b;�_�F�����/���|�����_�(ȟ�)bSː��F����S]f�dj���9^\=��9xT\e�I,�9����`�S�"����3�A�MEo[p͕W���`Ha�{�0�>��g�a�A|18�|��d���þ�#Q�-|�?��o|k�dr����߃!���-��<��y���&#9&�JX��Kစt3�Y�6Ym�V�����	1�|?���F_^}bw���
'�P#�.P�ʶ0ϥ}�&A��"\��&p�P� [F)�?�O�#�8������?�'�"T��*}�����}�pW·�~���q��q@��cc�#/�q��^6a:�Ǎ�"k�Zke��3��P'��7����� ����-My�e4!ۜ�-���㶚�J���G��l��Tۋ��tM���FAF�HE�����3=;z�3��5��y��>��@�f����'F�1�XD����H��䭧_��_�?��J�Պ����嬍<Q�"MhY�r��W�S�1�Iɹ0����Jv�*%'��їdh/|���'�����M��2UW/�����5�������:ǸW�e�:s�@�XC~��A�vO���IZ>[�bD|�^����sY�s���O0��0]U?�)ـG��?����@�i@=�$�S��G����I��vg�\��F���H�A�Wgoլ���}�;�����8�ѩᦦ�u"li<#�����nx�xhh�N�D�)�'zw?+8HP+ڷ (��j��c��fּ��!~�1�AXO�ӟ�9�}��?@��s�2 Ɔ>������!��b�$�-%��W����'^Kc���;��� ��}�n�-�>��$Ã �5���|�C�0��F������'��?C�̽j�yi����"������8�T�����Pp'�@�Vr�k^'l	^� £) v�}����{-2�A��l�J]�_.
t�q@m��t2�����G�#~_��z�s�p� �u�*�a}J��@��>I� %.�e��8n*�Ay���E�
G�gT�����_X�6� ���D~��I]�q�h����G�w�Ɏ�#V�MH�nn=<��0���c/�1YQ���LOFR�EyZ�"�	��� �5�}�����&?��?g_���_�g.�� �� y�*�`<c��չ�ZG��������TPǯ�S���ۿ�����|���0���` �>�x�s����5@*a{�i��p0O�k���&<atu2v.N	�i���� р�� %ID�D����_
sP���_-*W��>/+���clC5�w����Y��#�R��k��
v���/�Ó�?��Χ���,(�6���a��?k���;�_,�B;Z��r���U��.]a�S�z�����M�-�3~��o�� �V 1 ����Ib�о���_��e�.9�B	�f��B�����JBxW�������A��T���k:y���U�����ఞg�a�������9�s��/�q�����l=`�?yo�0|�}3��f��k�A�m{�%�y2d<��$�/����G��p8� AZ0���!3������gB�5Ʉ�r.XI�F��<��^�@��W~'�L�=����r �!����.j�v����4��v��QLМ��]䠱�~Z���~L� <���2��01��2�p�#!u�� ���T�M���K�.&e��}PJ9m�8�ހ���'�+�짃���>:��.s#���o��e���[�®)��s�1KG�8^�ܰ܁=_�r�������Λ���[
Q��:% >�f|�^M��h|�͘����6���b�!9A��j�I�0�����p�Y\p8F�>G:z��|澹|t�_޳����n{�����>�^��g'Xt<~�������M	�k+��z� B��ωt��?7�}��ѡ�#�T���G���$| ����3a�PEK�0@�l�憶?����g���2�p��g3���W�z2JO1�d���:�%���_\d���b�X`��-�zb/���e���
�}\/�W��	_Xߜ���$%����%?s g��2��sN��;M-a�= �)�v?�뎤��g���#+s��ے(����D�@��EA�����(�̿�1M�~�	�>��Q'S�q��.E'�!.R�v�ʪ�W:���y�7<e�n�R�Ur��r>)C��hC${bzW��pd�����1 �et~��r�?W1�u1���a�c�r�������G�6x���5/�5�s�2}\�M���z¦?��%�?Y|~��z?X�#]�|K�� B���^�1 ����e�G��<�����\���G�#"r9�j��2;X y��Ga1���It�����a��,0HO���/,<���a�}�/�hM�Y�?ۉ?b�pB"=�[���9�#����`�~|���m@��@D���H������ �?ư���N
�$^0�R��ڨ��ǃ-����2r��xo�,xI��*�z�,c3�����W�8���q7��/j�@�G˔�?�+��֏��p���?/��,sG/�ƌ���A�у�)��m�`N��\ύ�Ӄ�r��4�Ř�g*�ArϨ�Cy+�P��eKt~������s������ xDOq�0�Ú�������� ~s�����#��L4�?y��'�\X�fhTK����v���u}�����3$�s1}��U!:>;�NL�����G�ʰ�u����J�D���i�,/ȚU�0�����y���c
���L�e�_~;��9�V�Ӎ���1l�C��>���+�E��������F@ӈ��9=�E��8`�K��M�y"�ʖ���i0����Ux�&:Oh��H�eU�L���o�F�/y⤱?U��L���}sx;B�Y|h�\�O�FY7/Xu���t��$��(�ʷ��Ѽ��n$:��8P��O����K�d'YA�c���T/�W�x�����"~G�9��s���3Z���� Ş�g=7��}���	�,g�Ü��G�8��g?�s?n:zˌT8�s��M{�w����#~O,:*L�w4~��co��V��c%jo�R�-�W�5[{���Y+DK�򥨢b�H5J��Dk������y��s>��Ϲ�u�}��������P�'�����Zl\~�C�����	�{|�����/~��(�h��+�a� ��^<�\W��gλ�0Aa=���b�m��X��OThpc�[؛�*00�\���M]�WW��l,���p�3W��Pw����_�4�'�@AyLK/�zo�m����$�
�k`�C�Ve�P�����)���ޯ��Xli�3�?��5�����i����#n`���J~f��EDX�A�g���N����S�W��}v�~ךV$\i�:=Ln�����o�~Ͼ�n�Mj1����pО����S�I%I��$�T��� gê	��KF����;1�%M�R����S�]"�;ۨK|tm�o��֪����;��D�'��sA��~�|Җ�bif8��{�ye�B�|w�����$^����?���:��j^�έ���57�����L���5����H�� j��I"%U}dggʧ,�F,G�4{
�QXtd���Aپ�I�9Ny*��4.��,H�L(�q�{�C��3�D*�|w�M�:"� ���B�k4��t�$L/�?J�չz0�o�A�k�(})��=�� g<.G�(TV�tc{���`����'�S,l�x���xyu'�u��`�y������ UŜ�%��_Z}։��x�)�v��̃%�]/о7����ot�1���F�s�&v~)�GWE��,����a���R���շ��V��P�up�'*'v\$�
��kۥg.*(BeQp���Ý���=���h���A�����k_	��,K��Q]���3�p����ޟ��2s�|��uwY���GO6�ԐN� }������v�v�S�u����]k$S��V%����s9�u���?;!�����{5g��&�Q�擄��[ه���~�o�P�$��mu���>r���w|�*���[��樺� �Qm�%�j�U���E�����ԺΥ=��;}T%}�� Â���:�5.�lW��>�J��'��P�������E�_���.oDD	T��9�a;�W�p����(�C�]�o~*�g�n=����{��o����˞��m�����
��x��h�Q���˂��i�����N�txnT�/�u���u��U9��M<҉N#xp�.g�����/`�}�� ����yw����OB��`�Df<���G�cy����\w�r�u#��=͕c���$0Ŗ��g������AXS#�P[IvnT���CG��>vtZ4O����x�����X��sZe�%��0��C|#��Lw����K�˽�?Җڻ�B>��C5�1���	j��(�li�����5D/B.%��]u0��Y������ӆ�cDے�rx��ԆTF������e,w���Y#�{k���̷&�.��2sC���ޙ�0��gg��!Nq�����=DxeyQ�!�%��m:&C�יˏ�E>,. ��x$����θ~Z��[��� ǲ@AR~����e"�I��.Q�}��P�ߦԚlh^��^V�&5,0��D�)<�e��bh���H���eZ_�]�}��ܚQĊĬ��6	�}a̦
L~���n�\�{���q��W�ҲҾ:��:~w�G�����L-��W�U~�"3��v��ز?��o�ٹyߋ���0�'#��j$`�Q<�x��?��2��k�����|��ɓ%z�7�@Ȯ�N�L��Bh��@�,+�.\�*�� ��,�7�w����2ny5=n�XsF�OC-���������{>E6݌�����f����E�!�-\CSx��*�`:)e�c�����Z��|B�@ٳ����Q����1m�Eo�vB0��:a.��\��ׅ�c�l���[��]�p���&��Y�f����r9�$����O呉������[�|ѱ�y��4ȃ/=n~6[I@�p�����
�b@]n#��*��h�"r¦|7=�YΌ�+�Ix��(�S�ٺ��H.;����M��k[���l}��kd���������^		��w�܄k:邽>�(�m���7͜���k�.	���ΐ8���L��2Fo�Ԅ6�D����C�lW!��Dv�b��K���
��[�8֢>��-��S��Z����()J�n��ձ���e�}"Q	����H�V^�71��;K��Y�l�����k'��4egz;���c�S�l�	�X\*:^���`df.#��@d񷵌_��[�xGcE�u�G��t�ƈ4J��$-��À���|t�>�C�ܚ�52"�JG@�;w���-W�t؏�Gq�{�Fˆl�gM�:08U�V�S9�o���,
��3G=�#-�Մ�˃�^�8O�M�q=.<LڂD����.���{D4����6��̭Q�E�s���.?�%z(�c%�������ǡ���t{��k�g8�3�Q4/���4��hg+�n)���T��T��@w�K��D֯��.R�ɫxF	���s�}lΉ�c��̣{:v./l)A|��	i9��"����\�_�ŉw#�����Ր�����L���0BUݙ�$�+����o��_�8��a���-̯\�ԭ�<�6	bkRɱh�����䣀�+y��h�HZmy'l�R�����-D�O\t�dEt�:ՕN�4V�V���bF�w�M����3ҁ��yf��7ڿ3m��z/��v�� ���S�Zqm�^n�$�m��\lLT�����;&` ��v�������3@4�G��^�r]�I^V�����"V'�憼���K����V1���w���s�����
1�F�e�+C���`���O��f�26J6/���/9)����[r`�E� ��{?�^	}���G�C���<����f�9Wm��Rs �����c�4<�>�h�5C3�*�)������K����e"Fq���4�އ�1���O�J}�<[�Ҧ���ˁ�{���eSr�.��3>E3�ք�k{2!}�{�����d�7_�Jm�Gږ�D�%q���]v�2""��W��GN8B�c�@(�e�R�2Y�7E/�a�g��߁���EpN��Nn�Moc�&[[V$�@-�����L3�k��_���^w+��O��������]	�Z�	{_˖�S����h�`ޗ�;emJ���)ƻ��G�/��<�٧}v�`�d�gR\�ӎ� ��z
��U���ӵK��OKZ���=]>aq���}�us�'Q���8j���Z����=��{���
�"��9�siJ�u�3�׮R
rw��P9����W\�dBS3!��P�^qk���+ NUi	����l�I����C�1�[���@���?S��t釭l�����]�#��9D7��Z�A���ٻʉ�6��ΆT�B?"T�|m�1�I����%�M���L�^��}Y������,v1��ݬ��jM�	[gh�m?[��
w��@�4+n�
��jz�ň�S��8)��n=0]����p?�+Hq��W4��[����-��v��5͖��_��lP��t"�Q�W �kvs8͐�PG�^M��<5���K�1��羫ަ��f=,o��n"��x���M<�z�m� q�v���W��29�8"u�AۙDnH	}G�Z�헯�zL$��8��~G���u$B=�'-�Xu`ϊW�P����,׾�T����]�'�yyW����
V�P]�������qٿ�˂RN�18R�$	]�%�j��(,J��مMG����������`���Ɓ�b�VTʳ�!�s��� zr7H����<r>��zW�ޘ�"E�P���3~�CzmM�uW�}�E.W����!{�D3U;#�R��]�w��`phS_ē=?:�ҵ[��ݎ1ݿ�g��jAF"�}S�J���h�e��4t�.�S#�c��z:0�Tf�w�E1�xU-��?�;D���ӿU�_�g�.T��<��I��HG�U�(�x˕/>�[9��3�E����*j̏�� ��H���<��:,Pz~�E�|_�"�t0B��d1Ĩ��=�#Z]s��R/������a�����_$h��K���;k�h�СC�C��s��G����k���8��Vѐ��L�{<�.��~Fʗ7��A�H��J���~I�/��3�Խ���C���ڗ4���V�����ٞ�k���V8"g�pq�������z������v�GK�
Η��;訔�tIԺ&2QX�>�
�E�+Nj]�چ����^���&
E�����D��o����;#��l	�:q�>�IPi6ⲡ/�%��C�;B���v�>�趶��+�	mԏ׽ƪ�20O����
���]H�Q2�Uخ-[��)%�sk�CN�:)�na%���V�b-2�-�sۣ>�TP߲�Vh����E�Bmb�m	W���:>���% ���,�������Xi'=�N.�sQ:����B��'���hW�+�a���7I8����{jI4�GD�*��Ց�]H&C�OI��#��곴w��N=P��\/I%"���3�6�y�q��g�ƌ�����?�!c򯥕s$��E2.��4�������*(z|mB �z㳻%r���H˯i�c[}�����`�F�8�<
�A�5��^���xߝsA���k�^��������T{*[2��8p��MRJ��3�S�ۡ!�;q�5�}���2��A�#�]*���ܑ��֧�����Ix�}=����>��-�������19��o�`v���Ȭ�{=�GE��P��UB�n��s�!�o�"R��%���:��M�I�xG�{�/�W%w�x�D��=:����:������Y�L@��I���:��D��b6��V)j8Z�'l$�@jUn@�'U���]YJ������^��6����x�E
�|�]�D�b��]u$5��hU�(j��kf�k«�SL�|�\/Z�!��׌�8%�.��T�ʕ��BQ�@2_�����m�Ë~a?��GIY��3�9,Ch��#�]��W�
9R+�&�Wˏ���?b|M�zg��k1�^`f�w,E�F�ۅ�V�c�ϔx����F|6}E�S�H���K��w��n�ʵ�m�v�_='����I:���#�H���«Mt��C�U��aO�q���Aݧo��S7φB����"� �t6Ŷ�/����7�z�~����:%{�#�����ڣ�u�QE���8�����U��X��c�d������U�6�s�wi��Z�Eo.O�ѥ��L�fOm/�u�-*���/��ט��-��7N�����%����sk��E�@^*Z5�V5'>6R9����;�¿������J�4)Qm�ܾ���*EM��Q��K��j2�4���^�I��M���I5w�vw���{kЉ�Vj�=L�����|�����o�r���(]�?[{B��ɋ��f�_C0�vkh�KvL�x�	��:r{�2������f��J-_���z��)��% ����	q�,�<>�$�����[�j�,;,u,Z��4�m�,�ȡ.:���w������J�I����mu�v��/F��?�st�1|��X��w��a;8�g����q��d���T��m�[������d/ؤ�����bk�օ�Ҍ[!Y�9�D���кM2S>O-�݃�&w�W\'[)7���a}?��oX��T�����W��0����]¿�����ψ��<�֒�q}}�}_�hD�&��v��x�ϛu+<�v����8t�2�T�mC\�&d|��_OS�AQ�|��&(�A�irh���$�����F7/eL
I����@ވ_
z�5�$ǘx�m�<c%`�����G(��f|#��q��}��5����a�����Hÿ�+nќ�j+J�������h�Χ�5_��P��Xs�A���t�����g�,��E}|��GN,�-~�3Ez��	`��=�ֳs��7�[��W`]�� %�w�c��?��h��_~^�8&	����E�~�ۘ�#���f��D�b_���B���E��^����T)w�?�u��d�[M�>��G���Y��ӽ��7�D��ı 륆d�����r<�]�%	"���N�Ѯ"4o���`�#�ʬ?�ufc���Z�.K���c��g�����+Re���~uC�ޤ�-�\�����}�G�����{;��/n��^�E�1����ɥCԻ�kwDn�}|ڝ����c�ꚦ��F�]���|����>Ol;��rJ���p��2Is�ݏS*�Y}3t��y��qE���3�3Q��<�������:Ө����t�%!�;`M��G@�J���c����Wu�#�f����n�WE�F.ԝ�����B.�#`}ꁵ�;�Rڥ��|��̤�¦음�g
�L�+:b�h�j���:�����
M�FeZ:�Nc�ts\)1�1�&#Ei��{�"dkf:��ǖ����v<�"��������;4�Y�
 �x��z��g�~�)��!�n��V����4+�L����h��A�*���o�4��Ɔ����M��9���%�59���#%�͟
��ד���J��p�k�ym�E�h3s���Li��6&G�1gvx��pm{�7���ȹ���V�V<lh���)b{�>��1x�������	E)ݼ���ց��_�~h/����� �ˀHe���f9�D��n7�=I�2kd�vצ]!�0��#���wO3?��^Zn��.���-�y�I���]k̛�^}?�W���a���9;T=
\ǹ_� s���{%6)��l�JB�Җ��Ś(B���۴�Q !+�Q��e+�V�+�������~�l?`��0Sk7!�{<����ӧH�~���3꛶w��-�lo�*�����3����(���d����a���s�tM�)�9=����6�7�P��K���0X3|}�(�%���U���|X.P��竅��QI�2�Eخ͝��9ʹ J�K���W�{n.&���ۼ��U� [�cp��U�ԫi�au�F�{�l�D\,��(����q�ڤ�?j���|��E1ab���}�ޏ{�Q��4���ð4��+�Ҥ�=�:ё���oS�ǉ9[�������i?�^��)Ve�i	#V��n�a,\��o���{*����<�\�7�<Z��-�sV}�UlZ����%��B�ܡ�^6?ͪB�|��o��=^��7�睊��H����Jt�����V��Y�PG5%Y�SK,,vv&*��j�K��XK��H����/'�J��Z�~�f���]�V�k�ʍ��)�/��8EB�ˇ���M��zo�h�U_:ZK��6��JN������ O����k�}��!�	� fԊ�����u:���[��'ƙ����T!�e$�������Ʃ��ۈ� �p�[fD��59D�W2
�<+��z4���J�#���MєtUM7�ۜ��SL�p�q@��[c7��"i�fM�wLS�",O%8��Ar&�q�l�9v]���k2��(e��Zq���=1f�T�h60gJ���&�4i͵��g���_	o��RV>�6�S�����]����D��m%8N���hPYXv�7��2v���Uk����{��S�����5��3�<:ִE�9(����Pn�<�+ �֖�4O��nE^I���v9zL��b"��MqR:f��[��Gz4�Bi�sg�Ϧ
T��M$'ה
�L�W�jP�q�b3�O�x^�
���4�H֥�g@��K��pod�$P�t��Y��ݐ7�q�^�˧Oeh�E�;��z �q�%��Ͼ	P�3�YT��ep礥�9��S�˸ /�<�U�.X�$�����F|L)����@����ܼ���N�F���*�$��~/YQ�4�G�=����ʋx�þ�׹B׵m�.N�<�>�T�%mEW��'kv��ͨ���Ϯ G�"��f�6н�$µ$=OB��cv�=ȑ?��A4�w�t��a����ݖ;q�~޶@�&�yԺX	TBjW����Vp�W�d���5���� �& �+�K#Q�nGX�J��G��o��@���/2A�Q{�y��W Q���-%�;�4���yJ�8g��j���O�Ɍl���y��S1J����T� �Dr��^���.�Z(���,�®;D��z�Y������eϬk�:A�T9�4�[�R��x�o�2k����HK�i������;V�*˭Wd��CK-U��W��R�/��������fC��yR��0[BuL�|/-�_R�;��M����{���w�u�<�:E/Q�e]@,��ŵ޽K���%��q�dH7P�U���%�F�'&��%�A�v��K^ܜڢ����%W��%��36��8{%~O"2����h��gյ?[�]��6���� w�LE:�Ws�Y��Loo0�ܴ����ku݅�����Gŗy<V�q��WT�/�
W}@�p�n��g��+@O�	=�~GDE������؛�"	��6�[�<��.�0
k��s�eR���J�K��2Ja�(��%C� W���Py�T�pl�3��h�XP���7��W���U��L_}IKO<=tg���%-��rL��l)~���r�te0�'��$�}������j�=��}�'��Z�#��k�&d���@�y�wI���M�<J��s��(�a�WdJKm��l ���R,G�
����a4"��plҘ��y
��u�h_jz ��K�{Q��[�G�ώ+ F�����lV�_ୁ������;c�5�Q�������YY4D�Sp�/�o=�GO�GD)z�����UZ+�@2z��:��
r���-�K׼vT\��N��6�X�M�t\1̎�Jb��{�����̞pz
���3��o��t6�vw�C%�f;�޴�H��U�M��;�:c������
P��ƳE��e�s�	�u��&vX�hĝ��R��ΣZ�Cb��d��NW��^w�u[̗���L��F�J^����021�Jw�H`�;Q������NA�����{�!~�1\`�*�y��?�l]x���1O��l� 4����|��M:r�2P0�~��m�N���6�I9�$��:����6&���yo?9�r'��� �p�e\M����l��G\u.�:ҎEh�H���F\iIU�&��3���E��ֹ��F��;2�V�"���܋כ�e��R�L��M�fΝ�3�?_/����{R���F��R��*��)��{#�y���氩2�.�0�h�W�钸�dO��cN���g<�tr�(W	:H�Է-?����>P��K�������+�&ܜc�`f��.�o���V�M�����{@'���e�
�7OQ�3k�/1��Ƨ���D�@⫇�,��V���?�9(Q���-S�1<�פC&ǖ�Vf�T�v|:����;(�X�����aA��4��T�.�2zu7o'����_f�9�F���!
�gR���"�+��\9��k-HIVND,�Sf���J'1��\�aJt����lO�̅����D�֘�Aϼ�咑��@C�׳�,�ؘ��p!���.G�cG�6H�,٠�	V�?��1��t3y��;:ɮ(��*���wh��b:9�3�%�%G����2E��6�.nӽtI��^��$ �r�g���iڌ�v�������t���noOBB���1JP��%k�y��b�$��21&���}�Q����r�F�&5�.���{�
�t��ȳ���1뙿p�}ӟ��ׇ 5m[���C��X��5<q���L)|l/��)���,��}�*���ur����K%�xY�l����N���w�p�IsDM�@���@�q݁��򈛵�_�?�����!�x����h	>��xk�b��"��G)+�4;��u�e��'y��@�^�;8�(���E��������A��F��,���R�N�����_%؟x��Ѧ���{�(�Hʥ���)ه�/�_��ds�<�(ie�}����z��$��0�껿,�6��2`C�	S��b�9�m������?��������M0xڄ�yͯ�q�c�Z�!��v.⁄�tk�W ��3�(dL��϶}9���NvW��S3(_�Y�M�M)㿖2c�.L�q��ߌ�7xW�?���R�.t�ι�N�=V�Yc��R|�:ĵr�]'��VA�1%WF27��+���a���!ͥn�=֚��j��w��d���
���.��e�i�d��b� k�����FƍBQ{�#��7��s���j)T�u*��N�3sQ�ǁ�������H�(��2'��"��Ne��}_�J��`�� =��K�'�O�	�FK�b��Ǌ揇���5��ϣ}�6���;����l���1�2z$x�����v��|��.3�[�N:q��~���� �i�PbN�,C��/����Ӄ8��?ٷ�`���ƹA���_?���s�9��Z��k�)|W&R�H�7\o�B��b�{U�V���t` �R�1�f����-�r��imJ�7�9�yǔ��H�/̒?7k6@d���;�"֊��!�=��������isD>'�s|H@��jy��w*F1*���9j���^f2ĳ�r�<c0�Sb隋�?�RbR��8��Ę	��\g22���ҝ�5?�����c%�	^�Tn<_E��j&hr���1Q����6y[�BR�{~�F�'+����$I�]V_���φ#�~O7f7�rU�����=�j#��sZ�͘W�UP}��^���U4�a��s��ds*T�v��R[D|)f�}9����(2F�U�/�ٜ��G4��u��V����z�^�:4cY�R��:�t֤��r��S��U[m�Y��c'�����LI%�¢��h9T܅����ۚBqINe�p�7��!Nɠ���+��%X9$E]�E��YZ�M3[�4U�~V=�>���~���CQI�T}���� �Ps�bY�c=�?�䲙�hX[0���C�b����WM��r)��?���m�a���`�:@q�t\R4A�{ʟg�&�-tv�0�����S����e(��f�
P擬ற��z=-�U}�'����6�e��m\煫�A�]��e&]�=@3�y��t����G�"�@=4� G>�	�,dW,��o��?&��L�~��3j�?~��h�o�b-����Q�T;�Etw�`�P;7�t+A�Jѳ�8��O5�n�~ɰ?�̂$�l��W���� �.c�C���%^�G��@�x�b8V43�x�+�N�����T�[G�x��Gz�8d�|����R�/v��{���)��"*�y"bJ<�C0]7^*!��������c	��qVL%[f)�zÇuՃ��'������W���*��!>_�RB�g�x`�]�氡���͚@y�������gE��m�d��+�f�y�Y�t���}���P}C���l��+T�U��#2(:z�v�{ۤ`�k�*rLI��!?kf�i 茨Ʀ�ӵ�,@=g�-��5h��������<��_�l�ס����e]<xdR��3�6�Z\hF�O�*T�w��h'���XJ��I�a����f�FL��ْQ���ZP쉉LO��.�
{��%�!Z�oܙ�7_��@���.�.M�M��ė�]���S-Z����Uޯ���������&����l{�R�d�vzm
�v�
	��Թ��@�pϞ2c�^;�7򀡠$n�#ѕ������**���`�v� X{~Y�-C��C����	k�ZLo��mqBC�uƿ5 IJ|�X
B]������&X��_<�^pl����
T��AǙ�1P����м���Ŗ'�Eюx�V�(�HI��S�a� Z�k��J���6'F0؄<�Ȱk��|��?���7�6J��`��Rh�m����
��9�����K�M����X���(��.�%��4`@�')EV��ݧna<�4����}s
ΤqO�����8�NR�A����xB�N4T�z�	p�K���MD�GRÝ�
 �Ñ�X`P�,�������u�т0��>Z�Ԗ�����2�&'��2Cm��v�%+��<���`�w^�� ��;�u�7w�xb�6�cKׯI}zEǸ
���h�e�rB�"�R�^���V�o�Ӿ�~�չ �����M��6ptN�)�j���#G5h���C�w�^�ٖqՅ30`DO�h�Be�x4�*��%^�l������� ��](��~/���T���(�;��%!��G��E�"�`َ��Sz������@��Ҫ����<�o��Ue�<�[��u�p��[ܣg��Jm�~��g� �=oV�gꎿ�9�UHN7�����_�&�a~<��Sd���x��󛦥%oq�W����R���Y�05�WID����>��D�8�Y>G���d��	d��"�NA��7�a�(g\#G���"��6T[j�-�V�lx߷Y�_otϵ�.̰�t#%ި����)�-TV|,-,��(���%:"�����K�ōZTu8Ot\j��J�=��F�3�7�@���aI	wB|��Sϓ���虱q@@��[����$I��g���]�q(��Y�hp������@}s��_��.�TC���5�2�k�\�s�Q���	a��l���m���{�=�%�Wn^�a�j�C+R�-n�=6|M]7UF5[O��g�lXq�� ��$�1�סr��LN�m��F��4&�����0�֌�]�ա�Œ��De��~h�;�+���bQ�w�����8�)]�d/���YU"ߒ��������N�D��nS=5O&!W�s>�	�V2F������6���Æ��	Ț+�����ʔ���N�AB=i�Er�Z��~��z�`��<�~@��<;����%>�<�5{0Ǟl-�T����_��K\6gm����?��N=b'&N02F������7K�S��at
v�)��~�.[4#u3�V�&�P�X�O��м���썹�T�����X���i����M�Q��~`�����^��+���5��.��U�3����'wkq|)d��f���V�Lij{�${�X����g9��c��t���7�U���G�Ƕc^D�A���:gۦs�Y?�0ifr
g�m�y����V����}������F��J�̨���"§X�/�����ڮ��y��q���;e�Y;06?
XK�&��F���P'կ��Y!�1�A+q=��*�"$�D3;/��a��%��/:�BU&�]L$w�iۿ�#��@��`���IE�-faY�$��<=�҂A�ڭ�7�״�y�N3���aO2`���U��<=�`>	��q�WCg.��Cձ�(��6Ah�)�I:V~�v�v�
P���AD_����{�+��gg-}��� �@)M;ʯ��V�U�j;��H�<���BNF��-����G#�ē/��P�m�H���@ӡ�y�%-��mJҸ�����B�����D��>r�PS��<�,D]� ���W��-I��e�\�K��-Z)��C�5Ih]x��@��D\l�Q��ܨ=:¥��R͑� =�>��O��4!�X[B����T��z�U�6��Z�N��N��6m%!ԛo9U_e�F���G��U��&=�"W$��� f���ᦼ�&;sW��K�A0+,=��@�6��ߴ�3#W�$��
��<ۈ^.���K3$�6zU�
 G��9%� ��:� ��h�P�͡��Rg��W�
P��Q��������{� '��%�K_p���G_� �'�c�|N�>��.AE_b�� �ڿ�3�)���91n��=t�2[���c#*"*kc@?����o@��CenS����~�t�����,�{r���7j Sh�W�>��i$L93�_�4Գ��Q����W] �"1	���@�D�(%F�� א�{;�+�?���[�>��,Ɏ��k�.�	-���y���V�,{�bT��4D&k<V�q�f�sN�/(p�N��
�s�}y��$��U1>��O.U���pP���٠��2��e��,���@a��4i����=~T/�d�ˀ�m�o�*v�Zy���"��t�IQ�W�����{�^e��U�]�H)����m�8�%Yk�fP�~ǯ�zZʾ��*�AX"����H�;����
�r��O��avlc�/S��j�l�r��z����ˮ��=���M�6�w>f����8ے�`P��b࡬�Q١���@}J�r�[A)��u���M�KS
��V��H1��)�0�� �,s���t�L����L�%a2�b�G5< b<�ͥ�BSRxp5��5�Xj\��O�5x�+h�5��X��v���k��=� dz}�����IFo�N�y��VP]z��j� 
JjJ:Z*����@�.���w���C������nlþ�}��1NQ��kL���,�����A��<?�
�I��I7��	�, �;U��TZ��ߨQs���.�U���f^���.u��3��^��R�J��D7a�JP��_èu�F�Bԃ���l�RR��ǟ��S�w�,�*�fU7S����Z�s�]���;�Ǧ�W�T��z0
�t����>c��6��6�NHŀa������q��{���r���^5)���������w���a�����Y?�iM{aWb>/1 }���6�:%]�p�U�O���K�״��+�������|4;������|��
��s�tz��셕��A�������jQ�{�q"@9�/cl�.��#UF�~BaU؏;:���eC����X~��l�@��b��v�/�T�J6�6������rԦ�T^&���ٽ�Q9Ht�~�����n����d?�ț�	���1&�)`��u���7|K��Zo�F� K�{.��B�^_`���D_�I���m��'�����ƿ�y���*7��Y�4�p1��5---=-����@Ů�!�d�)��I����=�l��c����.b�Yz]c�2��7;T���\�j{Զ�0X�;+��� ��rڭ�{]��OW�i6L*_��;�ZՊK5�)���i�̆D%ꔡg����5�Q��*k"?ӣ��5f�矨��&�l������y�8���6�jP}a_��7�13xa��Ң2Up��AY����T�����rl�?��KG�����ҧ���)I�g��G���1F*��~������9�
�{s�>����N����c��	n|�a��@����>���5���Ғ\5�����k'm�u!f����Aς��]��cL%ʗ��}���o�{���_d�]������Q6��lnd�9�	P�`�˭.=�o��V0��-����7��li�7��^j{��!^��ak�����㢾,;� ����A ��e����S�xq����Z	��~t�W[���2�����O1��/^a���n��)���Lu\��K���_���j�WS��1ΦI=%t�l�߳! �ٌ�Ӿ|�Wt�,bR�϶1�Kt��� @g�ih��e�r<uSk��ޔ�Ę� ��Ĭ2?��{G�Ӭ���(�7׶�L�4?�J/���Hh�l�|Д)����9�%���:�S���,�Z���UҚy�h��hp��Z�ey4�?�x!���	0����z�����x�Z�яbu"T�ۑ�'Yqm}�/C�4gk��Aӆm^��;(��C)9d����~(S&��]�����a�M��Oų9w�mc�o�d�FA��b4���Q��]����o	�N�()Lb}�h���C/���v�cC,cڒo�o�!��ۑZ8+ELbF`?��J�YR|a'Y��(^�����Q�䖨J��-
?�}"�/�������_R�����X�=6�+��]Lߖo�Yg��#��F��;�k��jH��v���i������C��u�'�#o�h���G�'�9�I!J'�m~��ޮ/��*���k���$�|��J�����5������k�Kؑ�3�����q�S�:�� >~r��I�&'n~q]�=�z�� L�$G�����=]�譐�p:�k�����l�Twy��Дx8�K�ˬ2=�WU5�
g���7]����n��%sd�������~Ѽ��?��_pr#A>qj��S��O0}��!l&\B�2���%g�vcp�R�?Gs��7{�^ˊ$̸��� �=p�1Q�sˢ��,�bȆ�^��|�2�!c�w�>9�����_<��r͍`w����4�nB>��
�������*� �� +U��b���_FօB$�	X A�dL��6ɢ0#Q�Q�����Q���Эa
�%dǘ�YH>� ҌQ7$��(%4�M3*��V�1Px0��,�))Qb�h�B�*��&
�j�U���g���L+5�7�v�Nʖ�PMh���X��Ē��%'�U��6�%Z0$^1���9R-�<z�@�d��(]��v����gkɒ�&�3���ד;^L�y3���ד%�EЛ;^L(�����(u/��PK   ΄6Vv��0  �     jsons/user_defined.json��]o�6������~3w��Ҭ���bI�Z����v� ��Q�L�e�dd_ْ��z�{x�l�k\۵m�46/Jk�i��6�*�F����6m]�?���I�ڱ�;�|��ub&?[76K6�����/���p���y��iPJ���rR�2d��BM�c��T��8r��^�^l���7��]gMQov�vq�/2G|T��p\]�We^A����z��ϪպŰH1>��[T��!b�=۲�{�!�Wf�i
��>�T뢍�]��+����$�S�Q|�X�)��U��_ֺJRێX����8�x����j�χA>9�?�!��i�/�㧃|v���lx�y�����8���x�e�������}ʃ_w��h0c�RSն�O��&V��)�y�.1ڵ�׉�?���D�yW�����T3'�4KB�&$T` 4&g90! ��わ��O���4�B�`����dqD)5�FDR���|<��c�!��r<|�����tp6�w�N���v���Xx�k:8����fd��|B����reC?=�'r����D��<�ȡ���9���|"�~~��ܷ�:�~ݼZL6��׶tVf��.�lL5W,�INB&y,CE�M���39�x������ɔ8V<�[�œh����O�$'L��vRv
���IO�=Z��/�/�_�/�1�G0���$B�ٌ<?*AC�tj�����y���"cD�w!a��sL��"�|Ϸ�l[ ������ O(���ܧ�ܟ�Lp�����O�͠�Vp0�rv��F�Mข���O�M�W��\z5���+����FrǗ��-_����w '�9���]L�s"��
�I*B�Ε���Z�)�T��0��)P������	D���04�G�5��h;D����.n<
�/�!��Z��y8�^� n�t�����@'X\��﬒����M���U��n�s�|*�09�PRL*6	�UIh2&Lf���ɻ��c?��?Rɧ��|� <S�$QL9�i�C������>�>�PK
   ΄6V ��<�p  ��                  cirkitFile.jsonPK
   |��T��� �' /             �p  images/13cec52d-3863-489f-91e2-31075f0cbf82.jpgPK
   ��T`J�'�(  �)  /             �x images/1e039584-5af2-406d-af07-82deb6d77547.jpgPK
   
��TB��(�  /             �� images/31ebd35d-3137-4c9c-9389-844452b616c5.pngPK
   L��T���"d. -y /             � images/4b94d0a1-8bca-4ba2-81d1-ddf4f146611c.jpgPK
   �Tj$;�  T  /             �� images/55269798-4c36-498f-9f6d-2f3e7c8d88bb.jpgPK
   ��U���[B� B� /             � 	 images/b676df13-73e2-41ea-8e8a-dc46dce3d5cb.jpgPK
   ΄6Vv��0  �               ��
 jsons/user_defined.jsonPK      �  ��
   